module FFT32 
( 
input wire clk_20,clk_100, reset_all,
input wire signed [15:0] x0, x1, x2, x3, x4, x5, x6, x7, x8, x9, x10, x11, x12, x13, x14, 
x15, x16, x17, x18, x19, x20, x21, x22, x23, x24, x25, x26, x27, x28, x29, x30, x31,
output reg signed [15:0] out_real_0, out_real_1, out_real_2, out_real_3, out_real_4, out_real_5, out_real_6, 
out_real_7, out_real_8, out_real_9, out_real_10, out_real_11, out_real_12, out_real_13, out_real_14, out_real_15, 
out_real_16, out_real_17, out_real_18, out_real_19, out_real_20, out_real_21, out_real_22, out_real_23, out_real_24, out_real_25,
 out_real_26, out_real_27, out_real_28, out_real_29, out_real_30, out_real_31, 
output reg signed [15:0] out_imag_0, out_imag_1, out_imag_2, out_imag_3, out_imag_4, out_imag_5,
 out_imag_6, out_imag_7, out_imag_8, out_imag_9, out_imag_10, out_imag_11, out_imag_12, out_imag_13, out_imag_14, 
 out_imag_15, out_imag_16, out_imag_17, out_imag_18, out_imag_19, out_imag_20, out_imag_21, out_imag_22, out_imag_23,
 out_imag_24, out_imag_25, out_imag_26, out_imag_27, out_imag_28, out_imag_29, out_imag_30, out_imag_31

);
wire signed [15:0] w0_real=16'b0000000100000000 ;
wire signed [15:0] w0_imag=16'b0000000000000000 ;

wire signed [15:0] w1_real=16'b0000000011111011 ;
wire signed [15:0] w1_imag=16'b1111111111001111 ;

wire signed [15:0] w2_real=16'b0000000011101100 ;
wire signed [15:0] w2_imag=16'b1111111110011111 ;

wire signed [15:0] w3_real=16'b0000000011010100 ;
wire signed [15:0] w3_imag=16'b1111111101110010 ;

wire signed [15:0] w4_real=16'b0000000010110101 ;
wire signed [15:0] w4_imag=16'b1111111101001011 ;

wire signed [15:0] w5_real=16'b0000000010001110 ;
wire signed [15:0] w5_imag=16'b1111111100101100 ;

wire signed [15:0] w6_real=16'b0000000001100001 ;
wire signed [15:0] w6_imag=16'b1111111100010100 ;

wire signed [15:0] w7_real=16'b0000000000110001 ;
wire signed [15:0] w7_imag=16'b1111111100000101 ;

wire signed [15:0] w8_real=16'b0000000000000000 ;
wire signed [15:0] w8_imag=16'b1111111100000000 ;

wire signed [15:0] w9_real=16'b1111111111001111 ;
wire signed [15:0] w9_imag=16'b1111111100000101 ;

wire signed [15:0] w10_real=16'b1111111110011111 ;
wire signed [15:0] w10_imag=16'b1111111100010100 ;

wire signed [15:0] w11_real=16'b1111111101110010 ;
wire signed [15:0] w11_imag=16'b1111111100101100 ;

wire signed [15:0] w12_real=16'b1111111101001011 ;
wire signed [15:0] w12_imag=16'b1111111101001011 ;

wire signed [15:0] w13_real=16'b1111111100101100 ;
wire signed [15:0] w13_imag=16'b1111111101110010 ;

wire signed [15:0] w14_real=16'b1111111100010100 ;
wire signed [15:0] w14_imag=16'b1111111110011111 ;

wire signed [15:0] w15_real=16'b1111111100000101 ;
wire signed [15:0] w15_imag=16'b1111111111001111 ;

wire signed sload_s1 ,sload_s2, sload_s3, sload_s4, sload_s5;
wire signed aclr_s1, aclr_s2, aclr_s3, aclr_s4, aclr_s5;
wire signed [2:0] counter_out;
wire signed [15:0] stage1_in_real_0;
wire signed [15:0] stage1_in_imag_0;
wire signed [15:0] stage1_in_real_1;
wire signed [15:0] stage1_in_imag_1;
wire signed [15:0] stage1_in_real_2;
wire signed [15:0] stage1_in_imag_2;
wire signed [15:0] stage1_in_real_3;
wire signed [15:0] stage1_in_imag_3;
wire signed [15:0] stage1_in_real_4;
wire signed [15:0] stage1_in_imag_4;
wire signed [15:0] stage1_in_real_5;
wire signed [15:0] stage1_in_imag_5;
wire signed [15:0] stage1_in_real_6;
wire signed [15:0] stage1_in_imag_6;
wire signed [15:0] stage1_in_real_7;
wire signed [15:0] stage1_in_imag_7;
wire signed [15:0] stage1_in_real_8;
wire signed [15:0] stage1_in_imag_8;
wire signed [15:0] stage1_in_real_9;
wire signed [15:0] stage1_in_imag_9;
wire signed [15:0] stage1_in_real_10;
wire signed [15:0] stage1_in_imag_10;
wire signed [15:0] stage1_in_real_11;
wire signed [15:0] stage1_in_imag_11;
wire signed [15:0] stage1_in_real_12;
wire signed [15:0] stage1_in_imag_12;
wire signed [15:0] stage1_in_real_13;
wire signed [15:0] stage1_in_imag_13;
wire signed [15:0] stage1_in_real_14;
wire signed [15:0] stage1_in_imag_14;
wire signed [15:0] stage1_in_real_15;
wire signed [15:0] stage1_in_imag_15;
wire signed [15:0] stage1_in_real_16;
wire signed [15:0] stage1_in_imag_16;
wire signed [15:0] stage1_in_real_17;
wire signed [15:0] stage1_in_imag_17;
wire signed [15:0] stage1_in_real_18;
wire signed [15:0] stage1_in_imag_18;
wire signed [15:0] stage1_in_real_19;
wire signed [15:0] stage1_in_imag_19;
wire signed [15:0] stage1_in_real_20;
wire signed [15:0] stage1_in_imag_20;
wire signed [15:0] stage1_in_real_21;
wire signed [15:0] stage1_in_imag_21;
wire signed [15:0] stage1_in_real_22;
wire signed [15:0] stage1_in_imag_22;
wire signed [15:0] stage1_in_real_23;
wire signed [15:0] stage1_in_imag_23;
wire signed [15:0] stage1_in_real_24;
wire signed [15:0] stage1_in_imag_24;
wire signed [15:0] stage1_in_real_25;
wire signed [15:0] stage1_in_imag_25;
wire signed [15:0] stage1_in_real_26;
wire signed [15:0] stage1_in_imag_26;
wire signed [15:0] stage1_in_real_27;
wire signed [15:0] stage1_in_imag_27;
wire signed [15:0] stage1_in_real_28;
wire signed [15:0] stage1_in_imag_28;
wire signed [15:0] stage1_in_real_29;
wire signed [15:0] stage1_in_imag_29;
wire signed [15:0] stage1_in_real_30;
wire signed [15:0] stage1_in_imag_30;
wire signed [15:0] stage1_in_real_31;
wire signed [15:0] stage1_in_imag_31;
wire signed [15:0] stage2_in_real_0;
wire signed [15:0] stage2_in_imag_0;
wire signed [15:0] stage2_in_real_1;
wire signed [15:0] stage2_in_imag_1;
wire signed [15:0] stage2_in_real_2;
wire signed [15:0] stage2_in_imag_2;
wire signed [15:0] stage2_in_real_3;
wire signed [15:0] stage2_in_imag_3;
wire signed [15:0] stage2_in_real_4;
wire signed [15:0] stage2_in_imag_4;
wire signed [15:0] stage2_in_real_5;
wire signed [15:0] stage2_in_imag_5;
wire signed [15:0] stage2_in_real_6;
wire signed [15:0] stage2_in_imag_6;
wire signed [15:0] stage2_in_real_7;
wire signed [15:0] stage2_in_imag_7;
wire signed [15:0] stage2_in_real_8;
wire signed [15:0] stage2_in_imag_8;
wire signed [15:0] stage2_in_real_9;
wire signed [15:0] stage2_in_imag_9;
wire signed [15:0] stage2_in_real_10;
wire signed [15:0] stage2_in_imag_10;
wire signed [15:0] stage2_in_real_11;
wire signed [15:0] stage2_in_imag_11;
wire signed [15:0] stage2_in_real_12;
wire signed [15:0] stage2_in_imag_12;
wire signed [15:0] stage2_in_real_13;
wire signed [15:0] stage2_in_imag_13;
wire signed [15:0] stage2_in_real_14;
wire signed [15:0] stage2_in_imag_14;
wire signed [15:0] stage2_in_real_15;
wire signed [15:0] stage2_in_imag_15;
wire signed [15:0] stage2_in_real_16;
wire signed [15:0] stage2_in_imag_16;
wire signed [15:0] stage2_in_real_17;
wire signed [15:0] stage2_in_imag_17;
wire signed [15:0] stage2_in_real_18;
wire signed [15:0] stage2_in_imag_18;
wire signed [15:0] stage2_in_real_19;
wire signed [15:0] stage2_in_imag_19;
wire signed [15:0] stage2_in_real_20;
wire signed [15:0] stage2_in_imag_20;
wire signed [15:0] stage2_in_real_21;
wire signed [15:0] stage2_in_imag_21;
wire signed [15:0] stage2_in_real_22;
wire signed [15:0] stage2_in_imag_22;
wire signed [15:0] stage2_in_real_23;
wire signed [15:0] stage2_in_imag_23;
wire signed [15:0] stage2_in_real_24;
wire signed [15:0] stage2_in_imag_24;
wire signed [15:0] stage2_in_real_25;
wire signed [15:0] stage2_in_imag_25;
wire signed [15:0] stage2_in_real_26;
wire signed [15:0] stage2_in_imag_26;
wire signed [15:0] stage2_in_real_27;
wire signed [15:0] stage2_in_imag_27;
wire signed [15:0] stage2_in_real_28;
wire signed [15:0] stage2_in_imag_28;
wire signed [15:0] stage2_in_real_29;
wire signed [15:0] stage2_in_imag_29;
wire signed [15:0] stage2_in_real_30;
wire signed [15:0] stage2_in_imag_30;
wire signed [15:0] stage2_in_real_31;
wire signed [15:0] stage2_in_imag_31;
wire signed [15:0] stage3_in_real_0;
wire signed [15:0] stage3_in_imag_0;
wire signed [15:0] stage3_in_real_1;
wire signed [15:0] stage3_in_imag_1;
wire signed [15:0] stage3_in_real_2;
wire signed [15:0] stage3_in_imag_2;
wire signed [15:0] stage3_in_real_3;
wire signed [15:0] stage3_in_imag_3;
wire signed [15:0] stage3_in_real_4;
wire signed [15:0] stage3_in_imag_4;
wire signed [15:0] stage3_in_real_5;
wire signed [15:0] stage3_in_imag_5;
wire signed [15:0] stage3_in_real_6;
wire signed [15:0] stage3_in_imag_6;
wire signed [15:0] stage3_in_real_7;
wire signed [15:0] stage3_in_imag_7;
wire signed [15:0] stage3_in_real_8;
wire signed [15:0] stage3_in_imag_8;
wire signed [15:0] stage3_in_real_9;
wire signed [15:0] stage3_in_imag_9;
wire signed [15:0] stage3_in_real_10;
wire signed [15:0] stage3_in_imag_10;
wire signed [15:0] stage3_in_real_11;
wire signed [15:0] stage3_in_imag_11;
wire signed [15:0] stage3_in_real_12;
wire signed [15:0] stage3_in_imag_12;
wire signed [15:0] stage3_in_real_13;
wire signed [15:0] stage3_in_imag_13;
wire signed [15:0] stage3_in_real_14;
wire signed [15:0] stage3_in_imag_14;
wire signed [15:0] stage3_in_real_15;
wire signed [15:0] stage3_in_imag_15;
wire signed [15:0] stage3_in_real_16;
wire signed [15:0] stage3_in_imag_16;
wire signed [15:0] stage3_in_real_17;
wire signed [15:0] stage3_in_imag_17;
wire signed [15:0] stage3_in_real_18;
wire signed [15:0] stage3_in_imag_18;
wire signed [15:0] stage3_in_real_19;
wire signed [15:0] stage3_in_imag_19;
wire signed [15:0] stage3_in_real_20;
wire signed [15:0] stage3_in_imag_20;
wire signed [15:0] stage3_in_real_21;
wire signed [15:0] stage3_in_imag_21;
wire signed [15:0] stage3_in_real_22;
wire signed [15:0] stage3_in_imag_22;
wire signed [15:0] stage3_in_real_23;
wire signed [15:0] stage3_in_imag_23;
wire signed [15:0] stage3_in_real_24;
wire signed [15:0] stage3_in_imag_24;
wire signed [15:0] stage3_in_real_25;
wire signed [15:0] stage3_in_imag_25;
wire signed [15:0] stage3_in_real_26;
wire signed [15:0] stage3_in_imag_26;
wire signed [15:0] stage3_in_real_27;
wire signed [15:0] stage3_in_imag_27;
wire signed [15:0] stage3_in_real_28;
wire signed [15:0] stage3_in_imag_28;
wire signed [15:0] stage3_in_real_29;
wire signed [15:0] stage3_in_imag_29;
wire signed [15:0] stage3_in_real_30;
wire signed [15:0] stage3_in_imag_30;
wire signed [15:0] stage3_in_real_31;
wire signed [15:0] stage3_in_imag_31;
wire signed [15:0] stage4_in_real_0;
wire signed [15:0] stage4_in_imag_0;
wire signed [15:0] stage4_in_real_1;
wire signed [15:0] stage4_in_imag_1;
wire signed [15:0] stage4_in_real_2;
wire signed [15:0] stage4_in_imag_2;
wire signed [15:0] stage4_in_real_3;
wire signed [15:0] stage4_in_imag_3;
wire signed [15:0] stage4_in_real_4;
wire signed [15:0] stage4_in_imag_4;
wire signed [15:0] stage4_in_real_5;
wire signed [15:0] stage4_in_imag_5;
wire signed [15:0] stage4_in_real_6;
wire signed [15:0] stage4_in_imag_6;
wire signed [15:0] stage4_in_real_7;
wire signed [15:0] stage4_in_imag_7;
wire signed [15:0] stage4_in_real_8;
wire signed [15:0] stage4_in_imag_8;
wire signed [15:0] stage4_in_real_9;
wire signed [15:0] stage4_in_imag_9;
wire signed [15:0] stage4_in_real_10;
wire signed [15:0] stage4_in_imag_10;
wire signed [15:0] stage4_in_real_11;
wire signed [15:0] stage4_in_imag_11;
wire signed [15:0] stage4_in_real_12;
wire signed [15:0] stage4_in_imag_12;
wire signed [15:0] stage4_in_real_13;
wire signed [15:0] stage4_in_imag_13;
wire signed [15:0] stage4_in_real_14;
wire signed [15:0] stage4_in_imag_14;
wire signed [15:0] stage4_in_real_15;
wire signed [15:0] stage4_in_imag_15;
wire signed [15:0] stage4_in_real_16;
wire signed [15:0] stage4_in_imag_16;
wire signed [15:0] stage4_in_real_17;
wire signed [15:0] stage4_in_imag_17;
wire signed [15:0] stage4_in_real_18;
wire signed [15:0] stage4_in_imag_18;
wire signed [15:0] stage4_in_real_19;
wire signed [15:0] stage4_in_imag_19;
wire signed [15:0] stage4_in_real_20;
wire signed [15:0] stage4_in_imag_20;
wire signed [15:0] stage4_in_real_21;
wire signed [15:0] stage4_in_imag_21;
wire signed [15:0] stage4_in_real_22;
wire signed [15:0] stage4_in_imag_22;
wire signed [15:0] stage4_in_real_23;
wire signed [15:0] stage4_in_imag_23;
wire signed [15:0] stage4_in_real_24;
wire signed [15:0] stage4_in_imag_24;
wire signed [15:0] stage4_in_real_25;
wire signed [15:0] stage4_in_imag_25;
wire signed [15:0] stage4_in_real_26;
wire signed [15:0] stage4_in_imag_26;
wire signed [15:0] stage4_in_real_27;
wire signed [15:0] stage4_in_imag_27;
wire signed [15:0] stage4_in_real_28;
wire signed [15:0] stage4_in_imag_28;
wire signed [15:0] stage4_in_real_29;
wire signed [15:0] stage4_in_imag_29;
wire signed [15:0] stage4_in_real_30;
wire signed [15:0] stage4_in_imag_30;
wire signed [15:0] stage4_in_real_31;
wire signed [15:0] stage4_in_imag_31;
wire signed [15:0] stage5_in_real_0;
wire signed [15:0] stage5_in_imag_0;
wire signed [15:0] stage5_in_real_1;
wire signed [15:0] stage5_in_imag_1;
wire signed [15:0] stage5_in_real_2;
wire signed [15:0] stage5_in_imag_2;
wire signed [15:0] stage5_in_real_3;
wire signed [15:0] stage5_in_imag_3;
wire signed [15:0] stage5_in_real_4;
wire signed [15:0] stage5_in_imag_4;
wire signed [15:0] stage5_in_real_5;
wire signed [15:0] stage5_in_imag_5;
wire signed [15:0] stage5_in_real_6;
wire signed [15:0] stage5_in_imag_6;
wire signed [15:0] stage5_in_real_7;
wire signed [15:0] stage5_in_imag_7;
wire signed [15:0] stage5_in_real_8;
wire signed [15:0] stage5_in_imag_8;
wire signed [15:0] stage5_in_real_9;
wire signed [15:0] stage5_in_imag_9;
wire signed [15:0] stage5_in_real_10;
wire signed [15:0] stage5_in_imag_10;
wire signed [15:0] stage5_in_real_11;
wire signed [15:0] stage5_in_imag_11;
wire signed [15:0] stage5_in_real_12;
wire signed [15:0] stage5_in_imag_12;
wire signed [15:0] stage5_in_real_13;
wire signed [15:0] stage5_in_imag_13;
wire signed [15:0] stage5_in_real_14;
wire signed [15:0] stage5_in_imag_14;
wire signed [15:0] stage5_in_real_15;
wire signed [15:0] stage5_in_imag_15;
wire signed [15:0] stage5_in_real_16;
wire signed [15:0] stage5_in_imag_16;
wire signed [15:0] stage5_in_real_17;
wire signed [15:0] stage5_in_imag_17;
wire signed [15:0] stage5_in_real_18;
wire signed [15:0] stage5_in_imag_18;
wire signed [15:0] stage5_in_real_19;
wire signed [15:0] stage5_in_imag_19;
wire signed [15:0] stage5_in_real_20;
wire signed [15:0] stage5_in_imag_20;
wire signed [15:0] stage5_in_real_21;
wire signed [15:0] stage5_in_imag_21;
wire signed [15:0] stage5_in_real_22;
wire signed [15:0] stage5_in_imag_22;
wire signed [15:0] stage5_in_real_23;
wire signed [15:0] stage5_in_imag_23;
wire signed [15:0] stage5_in_real_24;
wire signed [15:0] stage5_in_imag_24;
wire signed [15:0] stage5_in_real_25;
wire signed [15:0] stage5_in_imag_25;
wire signed [15:0] stage5_in_real_26;
wire signed [15:0] stage5_in_imag_26;
wire signed [15:0] stage5_in_real_27;
wire signed [15:0] stage5_in_imag_27;
wire signed [15:0] stage5_in_real_28;
wire signed [15:0] stage5_in_imag_28;
wire signed [15:0] stage5_in_real_29;
wire signed [15:0] stage5_in_imag_29;
wire signed [15:0] stage5_in_real_30;
wire signed [15:0] stage5_in_imag_30;
wire signed [15:0] stage5_in_real_31;
wire signed [15:0] stage5_in_imag_31;



wire signed [15:0] stage1_out_real_0;
wire signed [15:0] stage1_out_imag_0;
wire signed [15:0] stage1_out_real_1;
wire signed [15:0] stage1_out_imag_1;
wire signed [15:0] stage1_out_real_2;
wire signed [15:0] stage1_out_imag_2;
wire signed [15:0] stage1_out_real_3;
wire signed [15:0] stage1_out_imag_3;
wire signed [15:0] stage1_out_real_4;
wire signed [15:0] stage1_out_imag_4;
wire signed [15:0] stage1_out_real_5;
wire signed [15:0] stage1_out_imag_5;
wire signed [15:0] stage1_out_real_6;
wire signed [15:0] stage1_out_imag_6;
wire signed [15:0] stage1_out_real_7;
wire signed [15:0] stage1_out_imag_7;
wire signed [15:0] stage1_out_real_8;
wire signed [15:0] stage1_out_imag_8;
wire signed [15:0] stage1_out_real_9;
wire signed [15:0] stage1_out_imag_9;
wire signed [15:0] stage1_out_real_10;
wire signed [15:0] stage1_out_imag_10;
wire signed [15:0] stage1_out_real_11;
wire signed [15:0] stage1_out_imag_11;
wire signed [15:0] stage1_out_real_12;
wire signed [15:0] stage1_out_imag_12;
wire signed [15:0] stage1_out_real_13;
wire signed [15:0] stage1_out_imag_13;
wire signed [15:0] stage1_out_real_14;
wire signed [15:0] stage1_out_imag_14;
wire signed [15:0] stage1_out_real_15;
wire signed [15:0] stage1_out_imag_15;
wire signed [15:0] stage1_out_real_16;
wire signed [15:0] stage1_out_imag_16;
wire signed [15:0] stage1_out_real_17;
wire signed [15:0] stage1_out_imag_17;
wire signed [15:0] stage1_out_real_18;
wire signed [15:0] stage1_out_imag_18;
wire signed [15:0] stage1_out_real_19;
wire signed [15:0] stage1_out_imag_19;
wire signed [15:0] stage1_out_real_20;
wire signed [15:0] stage1_out_imag_20;
wire signed [15:0] stage1_out_real_21;
wire signed [15:0] stage1_out_imag_21;
wire signed [15:0] stage1_out_real_22;
wire signed [15:0] stage1_out_imag_22;
wire signed [15:0] stage1_out_real_23;
wire signed [15:0] stage1_out_imag_23;
wire signed [15:0] stage1_out_real_24;
wire signed [15:0] stage1_out_imag_24;
wire signed [15:0] stage1_out_real_25;
wire signed [15:0] stage1_out_imag_25;
wire signed [15:0] stage1_out_real_26;
wire signed [15:0] stage1_out_imag_26;
wire signed [15:0] stage1_out_real_27;
wire signed [15:0] stage1_out_imag_27;
wire signed [15:0] stage1_out_real_28;
wire signed [15:0] stage1_out_imag_28;
wire signed [15:0] stage1_out_real_29;
wire signed [15:0] stage1_out_imag_29;
wire signed [15:0] stage1_out_real_30;
wire signed [15:0] stage1_out_imag_30;
wire signed [15:0] stage1_out_real_31;
wire signed [15:0] stage1_out_imag_31;
wire signed [15:0] stage2_out_real_0;
wire signed [15:0] stage2_out_imag_0;
wire signed [15:0] stage2_out_real_1;
wire signed [15:0] stage2_out_imag_1;
wire signed [15:0] stage2_out_real_2;
wire signed [15:0] stage2_out_imag_2;
wire signed [15:0] stage2_out_real_3;
wire signed [15:0] stage2_out_imag_3;
wire signed [15:0] stage2_out_real_4;
wire signed [15:0] stage2_out_imag_4;
wire signed [15:0] stage2_out_real_5;
wire signed [15:0] stage2_out_imag_5;
wire signed [15:0] stage2_out_real_6;
wire signed [15:0] stage2_out_imag_6;
wire signed [15:0] stage2_out_real_7;
wire signed [15:0] stage2_out_imag_7;
wire signed [15:0] stage2_out_real_8;
wire signed [15:0] stage2_out_imag_8;
wire signed [15:0] stage2_out_real_9;
wire signed [15:0] stage2_out_imag_9;
wire signed [15:0] stage2_out_real_10;
wire signed [15:0] stage2_out_imag_10;
wire signed [15:0] stage2_out_real_11;
wire signed [15:0] stage2_out_imag_11;
wire signed [15:0] stage2_out_real_12;
wire signed [15:0] stage2_out_imag_12;
wire signed [15:0] stage2_out_real_13;
wire signed [15:0] stage2_out_imag_13;
wire signed [15:0] stage2_out_real_14;
wire signed [15:0] stage2_out_imag_14;
wire signed [15:0] stage2_out_real_15;
wire signed [15:0] stage2_out_imag_15;
wire signed [15:0] stage2_out_real_16;
wire signed [15:0] stage2_out_imag_16;
wire signed [15:0] stage2_out_real_17;
wire signed [15:0] stage2_out_imag_17;
wire signed [15:0] stage2_out_real_18;
wire signed [15:0] stage2_out_imag_18;
wire signed [15:0] stage2_out_real_19;
wire signed [15:0] stage2_out_imag_19;
wire signed [15:0] stage2_out_real_20;
wire signed [15:0] stage2_out_imag_20;
wire signed [15:0] stage2_out_real_21;
wire signed [15:0] stage2_out_imag_21;
wire signed [15:0] stage2_out_real_22;
wire signed [15:0] stage2_out_imag_22;
wire signed [15:0] stage2_out_real_23;
wire signed [15:0] stage2_out_imag_23;
wire signed [15:0] stage2_out_real_24;
wire signed [15:0] stage2_out_imag_24;
wire signed [15:0] stage2_out_real_25;
wire signed [15:0] stage2_out_imag_25;
wire signed [15:0] stage2_out_real_26;
wire signed [15:0] stage2_out_imag_26;
wire signed [15:0] stage2_out_real_27;
wire signed [15:0] stage2_out_imag_27;
wire signed [15:0] stage2_out_real_28;
wire signed [15:0] stage2_out_imag_28;
wire signed [15:0] stage2_out_real_29;
wire signed [15:0] stage2_out_imag_29;
wire signed [15:0] stage2_out_real_30;
wire signed [15:0] stage2_out_imag_30;
wire signed [15:0] stage2_out_real_31;
wire signed [15:0] stage2_out_imag_31;
wire signed [15:0] stage3_out_real_0;
wire signed [15:0] stage3_out_imag_0;
wire signed [15:0] stage3_out_real_1;
wire signed [15:0] stage3_out_imag_1;
wire signed [15:0] stage3_out_real_2;
wire signed [15:0] stage3_out_imag_2;
wire signed [15:0] stage3_out_real_3;
wire signed [15:0] stage3_out_imag_3;
wire signed [15:0] stage3_out_real_4;
wire signed [15:0] stage3_out_imag_4;
wire signed [15:0] stage3_out_real_5;
wire signed [15:0] stage3_out_imag_5;
wire signed [15:0] stage3_out_real_6;
wire signed [15:0] stage3_out_imag_6;
wire signed [15:0] stage3_out_real_7;
wire signed [15:0] stage3_out_imag_7;
wire signed [15:0] stage3_out_real_8;
wire signed [15:0] stage3_out_imag_8;
wire signed [15:0] stage3_out_real_9;
wire signed [15:0] stage3_out_imag_9;
wire signed [15:0] stage3_out_real_10;
wire signed [15:0] stage3_out_imag_10;
wire signed [15:0] stage3_out_real_11;
wire signed [15:0] stage3_out_imag_11;
wire signed [15:0] stage3_out_real_12;
wire signed [15:0] stage3_out_imag_12;
wire signed [15:0] stage3_out_real_13;
wire signed [15:0] stage3_out_imag_13;
wire signed [15:0] stage3_out_real_14;
wire signed [15:0] stage3_out_imag_14;
wire signed [15:0] stage3_out_real_15;
wire signed [15:0] stage3_out_imag_15;
wire signed [15:0] stage3_out_real_16;
wire signed [15:0] stage3_out_imag_16;
wire signed [15:0] stage3_out_real_17;
wire signed [15:0] stage3_out_imag_17;
wire signed [15:0] stage3_out_real_18;
wire signed [15:0] stage3_out_imag_18;
wire signed [15:0] stage3_out_real_19;
wire signed [15:0] stage3_out_imag_19;
wire signed [15:0] stage3_out_real_20;
wire signed [15:0] stage3_out_imag_20;
wire signed [15:0] stage3_out_real_21;
wire signed [15:0] stage3_out_imag_21;
wire signed [15:0] stage3_out_real_22;
wire signed [15:0] stage3_out_imag_22;
wire signed [15:0] stage3_out_real_23;
wire signed [15:0] stage3_out_imag_23;
wire signed [15:0] stage3_out_real_24;
wire signed [15:0] stage3_out_imag_24;
wire signed [15:0] stage3_out_real_25;
wire signed [15:0] stage3_out_imag_25;
wire signed [15:0] stage3_out_real_26;
wire signed [15:0] stage3_out_imag_26;
wire signed [15:0] stage3_out_real_27;
wire signed [15:0] stage3_out_imag_27;
wire signed [15:0] stage3_out_real_28;
wire signed [15:0] stage3_out_imag_28;
wire signed [15:0] stage3_out_real_29;
wire signed [15:0] stage3_out_imag_29;
wire signed [15:0] stage3_out_real_30;
wire signed [15:0] stage3_out_imag_30;
wire signed [15:0] stage3_out_real_31;
wire signed [15:0] stage3_out_imag_31;
wire signed [15:0] stage4_out_real_0;
wire signed [15:0] stage4_out_imag_0;
wire signed [15:0] stage4_out_real_1;
wire signed [15:0] stage4_out_imag_1;
wire signed [15:0] stage4_out_real_2;
wire signed [15:0] stage4_out_imag_2;
wire signed [15:0] stage4_out_real_3;
wire signed [15:0] stage4_out_imag_3;
wire signed [15:0] stage4_out_real_4;
wire signed [15:0] stage4_out_imag_4;
wire signed [15:0] stage4_out_real_5;
wire signed [15:0] stage4_out_imag_5;
wire signed [15:0] stage4_out_real_6;
wire signed [15:0] stage4_out_imag_6;
wire signed [15:0] stage4_out_real_7;
wire signed [15:0] stage4_out_imag_7;
wire signed [15:0] stage4_out_real_8;
wire signed [15:0] stage4_out_imag_8;
wire signed [15:0] stage4_out_real_9;
wire signed [15:0] stage4_out_imag_9;
wire signed [15:0] stage4_out_real_10;
wire signed [15:0] stage4_out_imag_10;
wire signed [15:0] stage4_out_real_11;
wire signed [15:0] stage4_out_imag_11;
wire signed [15:0] stage4_out_real_12;
wire signed [15:0] stage4_out_imag_12;
wire signed [15:0] stage4_out_real_13;
wire signed [15:0] stage4_out_imag_13;
wire signed [15:0] stage4_out_real_14;
wire signed [15:0] stage4_out_imag_14;
wire signed [15:0] stage4_out_real_15;
wire signed [15:0] stage4_out_imag_15;
wire signed [15:0] stage4_out_real_16;
wire signed [15:0] stage4_out_imag_16;
wire signed [15:0] stage4_out_real_17;
wire signed [15:0] stage4_out_imag_17;
wire signed [15:0] stage4_out_real_18;
wire signed [15:0] stage4_out_imag_18;
wire signed [15:0] stage4_out_real_19;
wire signed [15:0] stage4_out_imag_19;
wire signed [15:0] stage4_out_real_20;
wire signed [15:0] stage4_out_imag_20;
wire signed [15:0] stage4_out_real_21;
wire signed [15:0] stage4_out_imag_21;
wire signed [15:0] stage4_out_real_22;
wire signed [15:0] stage4_out_imag_22;
wire signed [15:0] stage4_out_real_23;
wire signed [15:0] stage4_out_imag_23;
wire signed [15:0] stage4_out_real_24;
wire signed [15:0] stage4_out_imag_24;
wire signed [15:0] stage4_out_real_25;
wire signed [15:0] stage4_out_imag_25;
wire signed [15:0] stage4_out_real_26;
wire signed [15:0] stage4_out_imag_26;
wire signed [15:0] stage4_out_real_27;
wire signed [15:0] stage4_out_imag_27;
wire signed [15:0] stage4_out_real_28;
wire signed [15:0] stage4_out_imag_28;
wire signed [15:0] stage4_out_real_29;
wire signed [15:0] stage4_out_imag_29;
wire signed [15:0] stage4_out_real_30;
wire signed [15:0] stage4_out_imag_30;
wire signed [15:0] stage4_out_real_31;
wire signed [15:0] stage4_out_imag_31;
wire signed [15:0] stage5_out_real_0;
wire signed [15:0] stage5_out_imag_0;
wire signed [15:0] stage5_out_real_1;
wire signed [15:0] stage5_out_imag_1;
wire signed [15:0] stage5_out_real_2;
wire signed [15:0] stage5_out_imag_2;
wire signed [15:0] stage5_out_real_3;
wire signed [15:0] stage5_out_imag_3;
wire signed [15:0] stage5_out_real_4;
wire signed [15:0] stage5_out_imag_4;
wire signed [15:0] stage5_out_real_5;
wire signed [15:0] stage5_out_imag_5;
wire signed [15:0] stage5_out_real_6;
wire signed [15:0] stage5_out_imag_6;
wire signed [15:0] stage5_out_real_7;
wire signed [15:0] stage5_out_imag_7;
wire signed [15:0] stage5_out_real_8;
wire signed [15:0] stage5_out_imag_8;
wire signed [15:0] stage5_out_real_9;
wire signed [15:0] stage5_out_imag_9;
wire signed [15:0] stage5_out_real_10;
wire signed [15:0] stage5_out_imag_10;
wire signed [15:0] stage5_out_real_11;
wire signed [15:0] stage5_out_imag_11;
wire signed [15:0] stage5_out_real_12;
wire signed [15:0] stage5_out_imag_12;
wire signed [15:0] stage5_out_real_13;
wire signed [15:0] stage5_out_imag_13;
wire signed [15:0] stage5_out_real_14;
wire signed [15:0] stage5_out_imag_14;
wire signed [15:0] stage5_out_real_15;
wire signed [15:0] stage5_out_imag_15;
wire signed [15:0] stage5_out_real_16;
wire signed [15:0] stage5_out_imag_16;
wire signed [15:0] stage5_out_real_17;
wire signed [15:0] stage5_out_imag_17;
wire signed [15:0] stage5_out_real_18;
wire signed [15:0] stage5_out_imag_18;
wire signed [15:0] stage5_out_real_19;
wire signed [15:0] stage5_out_imag_19;
wire signed [15:0] stage5_out_real_20;
wire signed [15:0] stage5_out_imag_20;
wire signed [15:0] stage5_out_real_21;
wire signed [15:0] stage5_out_imag_21;
wire signed [15:0] stage5_out_real_22;
wire signed [15:0] stage5_out_imag_22;
wire signed [15:0] stage5_out_real_23;
wire signed [15:0] stage5_out_imag_23;
wire signed [15:0] stage5_out_real_24;
wire signed [15:0] stage5_out_imag_24;
wire signed [15:0] stage5_out_real_25;
wire signed [15:0] stage5_out_imag_25;
wire signed [15:0] stage5_out_real_26;
wire signed [15:0] stage5_out_imag_26;
wire signed [15:0] stage5_out_real_27;
wire signed [15:0] stage5_out_imag_27;
wire signed [15:0] stage5_out_real_28;
wire signed [15:0] stage5_out_imag_28;
wire signed [15:0] stage5_out_real_29;
wire signed [15:0] stage5_out_imag_29;
wire signed [15:0] stage5_out_real_30;
wire signed [15:0] stage5_out_imag_30;
wire signed [15:0] stage5_out_real_31;
wire signed [15:0] stage5_out_imag_31;


 controller_fsm conrtoller_i ( 
 .clk_100( clk_100 ),
 .clk_20( clk_20 ), .reset_all(reset_all),
.sload_s1(sload_s1) , .aclr_s1(aclr_s1) , 
.sload_s2(sload_s2) , .aclr_s2(aclr_s2) , 
.sload_s3(sload_s3) , .aclr_s3(aclr_s3) , 
.sload_s4(sload_s4) , .aclr_s4(aclr_s4) , 
.sload_s5(sload_s5) , .aclr_s5(aclr_s5) ,
.counter_out(  counter_out ));



Butterfly_C #(.data_width(16)) BF_1_0  (
.A_real( x0 ),.A_imag( 'd0), 
.B_real( x16 ), .B_imag( 'd0 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s1), .sload(sload_s1) 
,.select( counter_out[1:0]), .O_real(stage1_out_real_0  ), .O_imag( stage1_out_imag_0  ) );  

Butterfly_D #(.data_width(16)) BF_1_1  (
.A_real( x0 ),.A_imag( 'd0), 
.B_real( x16 ), .B_imag( 'd0 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s1), .sload(sload_s1) 
,.select( counter_out[1:0]), .O_real(stage1_out_real_1  ), .O_imag( stage1_out_imag_1  ) );  

/////////////////////////////////////////////////////////////////
Butterfly_C #(.data_width(16)) BF_1_2  (
.A_real( x1 ),.A_imag( 'd0), 
.B_real( x17 ), .B_imag( 'd0 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s1), .sload(sload_s1) 
,.select( counter_out[1:0]), .O_real(stage1_out_real_2  ), .O_imag( stage1_out_imag_2  ) );  

Butterfly_D #(.data_width(16)) BF_1_3  (
.A_real( x1 ),.A_imag( 'd0), 
.B_real( x17 ), .B_imag( 'd0 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s1), .sload(sload_s1) 
,.select( counter_out[1:0]), .O_real(stage1_out_real_3  ), .O_imag( stage1_out_imag_3  ) );  

/////////////////////////////////////////////////////////////////
Butterfly_C #(.data_width(16)) BF_1_4  (
.A_real( x2 ),.A_imag( 'd0), 
.B_real( x18 ), .B_imag( 'd0 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s1), .sload(sload_s1) 
,.select( counter_out[1:0]), .O_real(stage1_out_real_4  ), .O_imag( stage1_out_imag_4  ) );  

Butterfly_D #(.data_width(16)) BF_1_5  (
.A_real( x2 ),.A_imag( 'd0), 
.B_real( x18 ), .B_imag( 'd0 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s1), .sload(sload_s1) 
,.select( counter_out[1:0]), .O_real(stage1_out_real_5  ), .O_imag( stage1_out_imag_5  ) );  

/////////////////////////////////////////////////////////////////
Butterfly_C #(.data_width(16)) BF_1_6  (
.A_real( x3 ),.A_imag( 'd0), 
.B_real( x19 ), .B_imag( 'd0 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s1), .sload(sload_s1) 
,.select( counter_out[1:0]), .O_real(stage1_out_real_6  ), .O_imag( stage1_out_imag_6  ) );  

Butterfly_D #(.data_width(16)) BF_1_7  (
.A_real( x3 ),.A_imag( 'd0), 
.B_real( x19 ), .B_imag( 'd0 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s1), .sload(sload_s1) 
,.select( counter_out[1:0]), .O_real(stage1_out_real_7  ), .O_imag( stage1_out_imag_7  ) );  

/////////////////////////////////////////////////////////////////
Butterfly_C #(.data_width(16)) BF_1_8  (
.A_real( x4 ),.A_imag( 'd0), 
.B_real( x20 ), .B_imag( 'd0 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s1), .sload(sload_s1) 
,.select( counter_out[1:0]), .O_real(stage1_out_real_8  ), .O_imag( stage1_out_imag_8  ) );  

Butterfly_D #(.data_width(16)) BF_1_9  (
.A_real( x4 ),.A_imag( 'd0), 
.B_real( x20 ), .B_imag( 'd0 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s1), .sload(sload_s1) 
,.select( counter_out[1:0]), .O_real(stage1_out_real_9  ), .O_imag( stage1_out_imag_9  ) );  

/////////////////////////////////////////////////////////////////
Butterfly_C #(.data_width(16)) BF_1_10  (
.A_real( x5 ),.A_imag( 'd0), 
.B_real( x21 ), .B_imag( 'd0 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s1), .sload(sload_s1) 
,.select( counter_out[1:0]), .O_real(stage1_out_real_10  ), .O_imag( stage1_out_imag_10  ) );  

Butterfly_D #(.data_width(16)) BF_1_11  (
.A_real( x5 ),.A_imag( 'd0), 
.B_real( x21 ), .B_imag( 'd0 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s1), .sload(sload_s1) 
,.select( counter_out[1:0]), .O_real(stage1_out_real_11  ), .O_imag( stage1_out_imag_11  ) );  

/////////////////////////////////////////////////////////////////
Butterfly_C #(.data_width(16)) BF_1_12  (
.A_real( x6 ),.A_imag( 'd0), 
.B_real( x22 ), .B_imag( 'd0 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s1), .sload(sload_s1) 
,.select( counter_out[1:0]), .O_real(stage1_out_real_12  ), .O_imag( stage1_out_imag_12  ) );  

Butterfly_D #(.data_width(16)) BF_1_13  (
.A_real( x6 ),.A_imag( 'd0), 
.B_real( x22 ), .B_imag( 'd0 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s1), .sload(sload_s1) 
,.select( counter_out[1:0]), .O_real(stage1_out_real_13  ), .O_imag( stage1_out_imag_13  ) );  

/////////////////////////////////////////////////////////////////
Butterfly_C #(.data_width(16)) BF_1_14  (
.A_real( x7 ),.A_imag( 'd0), 
.B_real( x23 ), .B_imag( 'd0 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s1), .sload(sload_s1) 
,.select( counter_out[1:0]), .O_real(stage1_out_real_14  ), .O_imag( stage1_out_imag_14  ) );  

Butterfly_D #(.data_width(16)) BF_1_15  (
.A_real( x7 ),.A_imag( 'd0), 
.B_real( x23 ), .B_imag( 'd0 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s1), .sload(sload_s1) 
,.select( counter_out[1:0]), .O_real(stage1_out_real_15  ), .O_imag( stage1_out_imag_15  ) );  

/////////////////////////////////////////////////////////////////
Butterfly_C #(.data_width(16)) BF_1_16  (
.A_real( x8 ),.A_imag( 'd0), 
.B_real( x24 ), .B_imag( 'd0 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s1), .sload(sload_s1) 
,.select( counter_out[1:0]), .O_real(stage1_out_real_16  ), .O_imag( stage1_out_imag_16  ) );  

Butterfly_D #(.data_width(16)) BF_1_17  (
.A_real( x8 ),.A_imag( 'd0), 
.B_real( x24 ), .B_imag( 'd0 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s1), .sload(sload_s1) 
,.select( counter_out[1:0]), .O_real(stage1_out_real_17  ), .O_imag( stage1_out_imag_17  ) );  

/////////////////////////////////////////////////////////////////
Butterfly_C #(.data_width(16)) BF_1_18  (
.A_real( x9 ),.A_imag( 'd0), 
.B_real( x25 ), .B_imag( 'd0 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s1), .sload(sload_s1) 
,.select( counter_out[1:0]), .O_real(stage1_out_real_18  ), .O_imag( stage1_out_imag_18  ) );  

Butterfly_D #(.data_width(16)) BF_1_19  (
.A_real( x9 ),.A_imag( 'd0), 
.B_real( x25 ), .B_imag( 'd0 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s1), .sload(sload_s1) 
,.select( counter_out[1:0]), .O_real(stage1_out_real_19  ), .O_imag( stage1_out_imag_19  ) );  

/////////////////////////////////////////////////////////////////
Butterfly_C #(.data_width(16)) BF_1_20  (
.A_real( x10 ),.A_imag( 'd0), 
.B_real( x26 ), .B_imag( 'd0 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s1), .sload(sload_s1) 
,.select( counter_out[1:0]), .O_real(stage1_out_real_20  ), .O_imag( stage1_out_imag_20  ) );  

Butterfly_D #(.data_width(16)) BF_1_21  (
.A_real( x10 ),.A_imag( 'd0), 
.B_real( x26 ), .B_imag( 'd0 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s1), .sload(sload_s1) 
,.select( counter_out[1:0]), .O_real(stage1_out_real_21  ), .O_imag( stage1_out_imag_21  ) );  

/////////////////////////////////////////////////////////////////
Butterfly_C #(.data_width(16)) BF_1_22  (
.A_real( x11 ),.A_imag( 'd0), 
.B_real( x27 ), .B_imag( 'd0 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s1), .sload(sload_s1) 
,.select( counter_out[1:0]), .O_real(stage1_out_real_22  ), .O_imag( stage1_out_imag_22  ) );  

Butterfly_D #(.data_width(16)) BF_1_23  (
.A_real( x11 ),.A_imag( 'd0), 
.B_real( x27 ), .B_imag( 'd0 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s1), .sload(sload_s1) 
,.select( counter_out[1:0]), .O_real(stage1_out_real_23  ), .O_imag( stage1_out_imag_23  ) );  

/////////////////////////////////////////////////////////////////
Butterfly_C #(.data_width(16)) BF_1_24  (
.A_real( x12 ),.A_imag( 'd0), 
.B_real( x28 ), .B_imag( 'd0 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s1), .sload(sload_s1) 
,.select( counter_out[1:0]), .O_real(stage1_out_real_24  ), .O_imag( stage1_out_imag_24  ) );  

Butterfly_D #(.data_width(16)) BF_1_25  (
.A_real( x12 ),.A_imag( 'd0), 
.B_real( x28 ), .B_imag( 'd0 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s1), .sload(sload_s1) 
,.select( counter_out[1:0]), .O_real(stage1_out_real_25  ), .O_imag( stage1_out_imag_25  ) );  

/////////////////////////////////////////////////////////////////
Butterfly_C #(.data_width(16)) BF_1_26  (
.A_real( x13 ),.A_imag( 'd0), 
.B_real( x29 ), .B_imag( 'd0 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s1), .sload(sload_s1) 
,.select( counter_out[1:0]), .O_real(stage1_out_real_26  ), .O_imag( stage1_out_imag_26  ) );  

Butterfly_D #(.data_width(16)) BF_1_27  (
.A_real( x13 ),.A_imag( 'd0), 
.B_real( x29 ), .B_imag( 'd0 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s1), .sload(sload_s1) 
,.select( counter_out[1:0]), .O_real(stage1_out_real_27  ), .O_imag( stage1_out_imag_27  ) );  

/////////////////////////////////////////////////////////////////
Butterfly_C #(.data_width(16)) BF_1_28  (
.A_real( x14 ),.A_imag( 'd0), 
.B_real( x30 ), .B_imag( 'd0 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s1), .sload(sload_s1) 
,.select( counter_out[1:0]), .O_real(stage1_out_real_28  ), .O_imag( stage1_out_imag_28  ) );  

Butterfly_D #(.data_width(16)) BF_1_29  (
.A_real( x14 ),.A_imag( 'd0), 
.B_real( x30 ), .B_imag( 'd0 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s1), .sload(sload_s1) 
,.select( counter_out[1:0]), .O_real(stage1_out_real_29  ), .O_imag( stage1_out_imag_29  ) );  

/////////////////////////////////////////////////////////////////
Butterfly_C #(.data_width(16)) BF_1_30  (
.A_real( x15 ),.A_imag( 'd0), 
.B_real( x31 ), .B_imag( 'd0 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s1), .sload(sload_s1) 
,.select( counter_out[1:0]), .O_real(stage1_out_real_30  ), .O_imag( stage1_out_imag_30  ) );  

Butterfly_D #(.data_width(16)) BF_1_31  (
.A_real( x15 ),.A_imag( 'd0), 
.B_real( x31 ), .B_imag( 'd0 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s1), .sload(sload_s1) 
,.select( counter_out[1:0]), .O_real(stage1_out_real_31  ), .O_imag( stage1_out_imag_31  ) );  

/////////////////////////////////////////////////////////////////
Butterfly_C #(.data_width(16)) BF_2_0  (
.A_real(stage2_in_real_0),.A_imag( stage2_in_imag_0), 
.B_real( stage2_in_real_2 ), .B_imag(  stage2_in_imag_2 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s2), .sload(sload_s2) 
,.select( counter_out[1:0]), .O_real(stage2_out_real_0  ), .O_imag( stage2_out_imag_0  ) );  

Butterfly_C #(.data_width(16)) BF_2_1  (
.A_real(stage2_in_real_1),.A_imag( stage2_in_imag_1), 
.B_real(stage2_in_real_3 ), .B_imag( stage2_in_imag_3),
.W_real(  w8_real  ), .W_imag( w8_imag )
, .clk_MAC(clk_100), .aclr( aclr_s2), .sload(sload_s2) 
,.select( counter_out[1:0]), .O_real(stage2_out_real_1  ), .O_imag( stage2_out_imag_1  ) );  

Butterfly_D #(.data_width(16)) BF_2_2  (
.A_real(stage2_in_real_0),.A_imag( stage2_in_imag_0), 
.B_real(stage2_in_real_2 ), .B_imag(  stage2_in_imag_2 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s2), .sload(sload_s2) 
,.select( counter_out[1:0]), .O_real(stage2_out_real_2  ), .O_imag( stage2_out_imag_2  ) );  

Butterfly_D #(.data_width(16)) BF_2_3  (
.A_real(stage2_in_real_1),.A_imag( stage2_in_imag_1), 
.B_real( stage2_in_real_3 ), .B_imag(  stage2_in_imag_3 ),
.W_real(  w8_real  ), .W_imag( w8_imag )
, .clk_MAC(clk_100), .aclr( aclr_s2), .sload(sload_s2) 
,.select( counter_out[1:0]), .O_real(stage2_out_real_3  ), .O_imag( stage2_out_imag_3  ) );  

/////////////////////////////////////////////////////////////////
Butterfly_C #(.data_width(16)) BF_2_4  (
.A_real(stage2_in_real_4),.A_imag( stage2_in_imag_4), 
.B_real( stage2_in_real_6 ), .B_imag(  stage2_in_imag_6 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s2), .sload(sload_s2) 
,.select( counter_out[1:0]), .O_real(stage2_out_real_4  ), .O_imag( stage2_out_imag_4  ) );  

Butterfly_C #(.data_width(16)) BF_2_5  (
.A_real(stage2_in_real_5),.A_imag( stage2_in_imag_5), 
.B_real(stage2_in_real_7 ), .B_imag( stage2_in_imag_7),
.W_real(  w8_real  ), .W_imag( w8_imag )
, .clk_MAC(clk_100), .aclr( aclr_s2), .sload(sload_s2) 
,.select( counter_out[1:0]), .O_real(stage2_out_real_5  ), .O_imag( stage2_out_imag_5  ) );  

Butterfly_D #(.data_width(16)) BF_2_6  (
.A_real(stage2_in_real_4),.A_imag( stage2_in_imag_4), 
.B_real(stage2_in_real_6 ), .B_imag(  stage2_in_imag_6 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s2), .sload(sload_s2) 
,.select( counter_out[1:0]), .O_real(stage2_out_real_6  ), .O_imag( stage2_out_imag_6  ) );  

Butterfly_D #(.data_width(16)) BF_2_7  (
.A_real(stage2_in_real_5),.A_imag( stage2_in_imag_5), 
.B_real( stage2_in_real_7 ), .B_imag(  stage2_in_imag_7 ),
.W_real(  w8_real  ), .W_imag( w8_imag )
, .clk_MAC(clk_100), .aclr( aclr_s2), .sload(sload_s2) 
,.select( counter_out[1:0]), .O_real(stage2_out_real_7  ), .O_imag( stage2_out_imag_7  ) );  

/////////////////////////////////////////////////////////////////
Butterfly_C #(.data_width(16)) BF_2_8  (
.A_real(stage2_in_real_8),.A_imag( stage2_in_imag_8), 
.B_real( stage2_in_real_10 ), .B_imag(  stage2_in_imag_10 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s2), .sload(sload_s2) 
,.select( counter_out[1:0]), .O_real(stage2_out_real_8  ), .O_imag( stage2_out_imag_8  ) );  

Butterfly_C #(.data_width(16)) BF_2_9  (
.A_real(stage2_in_real_9),.A_imag( stage2_in_imag_9), 
.B_real(stage2_in_real_11 ), .B_imag( stage2_in_imag_11),
.W_real(  w8_real  ), .W_imag( w8_imag )
, .clk_MAC(clk_100), .aclr( aclr_s2), .sload(sload_s2) 
,.select( counter_out[1:0]), .O_real(stage2_out_real_9  ), .O_imag( stage2_out_imag_9  ) );  

Butterfly_D #(.data_width(16)) BF_2_10  (
.A_real(stage2_in_real_8),.A_imag( stage2_in_imag_8), 
.B_real(stage2_in_real_10 ), .B_imag(  stage2_in_imag_10 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s2), .sload(sload_s2) 
,.select( counter_out[1:0]), .O_real(stage2_out_real_10  ), .O_imag( stage2_out_imag_10  ) );  

Butterfly_D #(.data_width(16)) BF_2_11  (
.A_real(stage2_in_real_9),.A_imag( stage2_in_imag_9), 
.B_real( stage2_in_real_11 ), .B_imag(  stage2_in_imag_11 ),
.W_real(  w8_real  ), .W_imag( w8_imag )
, .clk_MAC(clk_100), .aclr( aclr_s2), .sload(sload_s2) 
,.select( counter_out[1:0]), .O_real(stage2_out_real_11  ), .O_imag( stage2_out_imag_11  ) );  

/////////////////////////////////////////////////////////////////
Butterfly_C #(.data_width(16)) BF_2_12  (
.A_real(stage2_in_real_12),.A_imag( stage2_in_imag_12), 
.B_real( stage2_in_real_14 ), .B_imag(  stage2_in_imag_14 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s2), .sload(sload_s2) 
,.select( counter_out[1:0]), .O_real(stage2_out_real_12  ), .O_imag( stage2_out_imag_12  ) );  

Butterfly_C #(.data_width(16)) BF_2_13  (
.A_real(stage2_in_real_13),.A_imag( stage2_in_imag_13), 
.B_real(stage2_in_real_15 ), .B_imag( stage2_in_imag_15),
.W_real(  w8_real  ), .W_imag( w8_imag )
, .clk_MAC(clk_100), .aclr( aclr_s2), .sload(sload_s2) 
,.select( counter_out[1:0]), .O_real(stage2_out_real_13  ), .O_imag( stage2_out_imag_13  ) );  

Butterfly_D #(.data_width(16)) BF_2_14  (
.A_real(stage2_in_real_12),.A_imag( stage2_in_imag_12), 
.B_real(stage2_in_real_14 ), .B_imag(  stage2_in_imag_14 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s2), .sload(sload_s2) 
,.select( counter_out[1:0]), .O_real(stage2_out_real_14  ), .O_imag( stage2_out_imag_14  ) );  

Butterfly_D #(.data_width(16)) BF_2_15  (
.A_real(stage2_in_real_13),.A_imag( stage2_in_imag_13), 
.B_real( stage2_in_real_15 ), .B_imag(  stage2_in_imag_15 ),
.W_real(  w8_real  ), .W_imag( w8_imag )
, .clk_MAC(clk_100), .aclr( aclr_s2), .sload(sload_s2) 
,.select( counter_out[1:0]), .O_real(stage2_out_real_15  ), .O_imag( stage2_out_imag_15  ) );  

/////////////////////////////////////////////////////////////////
Butterfly_C #(.data_width(16)) BF_2_16  (
.A_real(stage2_in_real_16),.A_imag( stage2_in_imag_16), 
.B_real( stage2_in_real_18 ), .B_imag(  stage2_in_imag_18 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s2), .sload(sload_s2) 
,.select( counter_out[1:0]), .O_real(stage2_out_real_16  ), .O_imag( stage2_out_imag_16  ) );  

Butterfly_C #(.data_width(16)) BF_2_17  (
.A_real(stage2_in_real_17),.A_imag( stage2_in_imag_17), 
.B_real(stage2_in_real_19 ), .B_imag( stage2_in_imag_19),
.W_real(  w8_real  ), .W_imag( w8_imag )
, .clk_MAC(clk_100), .aclr( aclr_s2), .sload(sload_s2) 
,.select( counter_out[1:0]), .O_real(stage2_out_real_17  ), .O_imag( stage2_out_imag_17  ) );  

Butterfly_D #(.data_width(16)) BF_2_18  (
.A_real(stage2_in_real_16),.A_imag( stage2_in_imag_16), 
.B_real(stage2_in_real_18 ), .B_imag(  stage2_in_imag_18 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s2), .sload(sload_s2) 
,.select( counter_out[1:0]), .O_real(stage2_out_real_18  ), .O_imag( stage2_out_imag_18  ) );  

Butterfly_D #(.data_width(16)) BF_2_19  (
.A_real(stage2_in_real_17),.A_imag( stage2_in_imag_17), 
.B_real( stage2_in_real_19 ), .B_imag(  stage2_in_imag_19 ),
.W_real(  w8_real  ), .W_imag( w8_imag )
, .clk_MAC(clk_100), .aclr( aclr_s2), .sload(sload_s2) 
,.select( counter_out[1:0]), .O_real(stage2_out_real_19  ), .O_imag( stage2_out_imag_19  ) );  

/////////////////////////////////////////////////////////////////
Butterfly_C #(.data_width(16)) BF_2_20  (
.A_real(stage2_in_real_20),.A_imag( stage2_in_imag_20), 
.B_real( stage2_in_real_22 ), .B_imag(  stage2_in_imag_22 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s2), .sload(sload_s2) 
,.select( counter_out[1:0]), .O_real(stage2_out_real_20  ), .O_imag( stage2_out_imag_20  ) );  

Butterfly_C #(.data_width(16)) BF_2_21  (
.A_real(stage2_in_real_21),.A_imag( stage2_in_imag_21), 
.B_real(stage2_in_real_23 ), .B_imag( stage2_in_imag_23),
.W_real(  w8_real  ), .W_imag( w8_imag )
, .clk_MAC(clk_100), .aclr( aclr_s2), .sload(sload_s2) 
,.select( counter_out[1:0]), .O_real(stage2_out_real_21  ), .O_imag( stage2_out_imag_21  ) );  

Butterfly_D #(.data_width(16)) BF_2_22  (
.A_real(stage2_in_real_20),.A_imag( stage2_in_imag_20), 
.B_real(stage2_in_real_22 ), .B_imag(  stage2_in_imag_22 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s2), .sload(sload_s2) 
,.select( counter_out[1:0]), .O_real(stage2_out_real_22  ), .O_imag( stage2_out_imag_22  ) );  

Butterfly_D #(.data_width(16)) BF_2_23  (
.A_real(stage2_in_real_21),.A_imag( stage2_in_imag_21), 
.B_real( stage2_in_real_23 ), .B_imag(  stage2_in_imag_23 ),
.W_real(  w8_real  ), .W_imag( w8_imag )
, .clk_MAC(clk_100), .aclr( aclr_s2), .sload(sload_s2) 
,.select( counter_out[1:0]), .O_real(stage2_out_real_23  ), .O_imag( stage2_out_imag_23  ) );  

/////////////////////////////////////////////////////////////////
Butterfly_C #(.data_width(16)) BF_2_24  (
.A_real(stage2_in_real_24),.A_imag( stage2_in_imag_24), 
.B_real( stage2_in_real_26 ), .B_imag(  stage2_in_imag_26 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s2), .sload(sload_s2) 
,.select( counter_out[1:0]), .O_real(stage2_out_real_24  ), .O_imag( stage2_out_imag_24  ) );  

Butterfly_C #(.data_width(16)) BF_2_25  (
.A_real(stage2_in_real_25),.A_imag( stage2_in_imag_25), 
.B_real(stage2_in_real_27 ), .B_imag( stage2_in_imag_27),
.W_real(  w8_real  ), .W_imag( w8_imag )
, .clk_MAC(clk_100), .aclr( aclr_s2), .sload(sload_s2) 
,.select( counter_out[1:0]), .O_real(stage2_out_real_25  ), .O_imag( stage2_out_imag_25  ) );  

Butterfly_D #(.data_width(16)) BF_2_26  (
.A_real(stage2_in_real_24),.A_imag( stage2_in_imag_24), 
.B_real(stage2_in_real_26 ), .B_imag(  stage2_in_imag_26 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s2), .sload(sload_s2) 
,.select( counter_out[1:0]), .O_real(stage2_out_real_26  ), .O_imag( stage2_out_imag_26  ) );  

Butterfly_D #(.data_width(16)) BF_2_27  (
.A_real(stage2_in_real_25),.A_imag( stage2_in_imag_25), 
.B_real( stage2_in_real_27 ), .B_imag(  stage2_in_imag_27 ),
.W_real(  w8_real  ), .W_imag( w8_imag )
, .clk_MAC(clk_100), .aclr( aclr_s2), .sload(sload_s2) 
,.select( counter_out[1:0]), .O_real(stage2_out_real_27  ), .O_imag( stage2_out_imag_27  ) );  

/////////////////////////////////////////////////////////////////
Butterfly_C #(.data_width(16)) BF_2_28  (
.A_real(stage2_in_real_28),.A_imag( stage2_in_imag_28), 
.B_real( stage2_in_real_30 ), .B_imag(  stage2_in_imag_30 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s2), .sload(sload_s2) 
,.select( counter_out[1:0]), .O_real(stage2_out_real_28  ), .O_imag( stage2_out_imag_28  ) );  

Butterfly_C #(.data_width(16)) BF_2_29  (
.A_real(stage2_in_real_29),.A_imag( stage2_in_imag_29), 
.B_real(stage2_in_real_31 ), .B_imag( stage2_in_imag_31),
.W_real(  w8_real  ), .W_imag( w8_imag )
, .clk_MAC(clk_100), .aclr( aclr_s2), .sload(sload_s2) 
,.select( counter_out[1:0]), .O_real(stage2_out_real_29  ), .O_imag( stage2_out_imag_29  ) );  

Butterfly_D #(.data_width(16)) BF_2_30  (
.A_real(stage2_in_real_28),.A_imag( stage2_in_imag_28), 
.B_real(stage2_in_real_30 ), .B_imag(  stage2_in_imag_30 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s2), .sload(sload_s2) 
,.select( counter_out[1:0]), .O_real(stage2_out_real_30  ), .O_imag( stage2_out_imag_30  ) );  

Butterfly_D #(.data_width(16)) BF_2_31  (
.A_real(stage2_in_real_29),.A_imag( stage2_in_imag_29), 
.B_real( stage2_in_real_31 ), .B_imag(  stage2_in_imag_31 ),
.W_real(  w8_real  ), .W_imag( w8_imag )
, .clk_MAC(clk_100), .aclr( aclr_s2), .sload(sload_s2) 
,.select( counter_out[1:0]), .O_real(stage2_out_real_31  ), .O_imag( stage2_out_imag_31  ) );  

/////////////////////////////////////////////////////////////////



Butterfly_C #(.data_width(16)) BF_3_0  (
.A_real( stage3_in_real_0 ),.A_imag( stage3_in_imag_0 ), 
.B_real( stage3_in_real_4 ), .B_imag( stage3_in_imag_4 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s3), .sload(sload_s3) 
,.select( counter_out[1:0]), .O_real(stage3_out_real_0  ), .O_imag( stage3_out_imag_0  ) );  

Butterfly_C #(.data_width(16)) BF_3_1  (
.A_real( stage3_in_real_1 ),.A_imag( stage3_in_imag_1 ), 
.B_real( stage3_in_real_5 ), .B_imag( stage3_in_imag_5 ),
.W_real(  w4_real  ), .W_imag( w4_imag )
, .clk_MAC(clk_100), .aclr( aclr_s3), .sload(sload_s3) 
,.select( counter_out[1:0]), .O_real(stage3_out_real_1  ), .O_imag( stage3_out_imag_1  ) );  

Butterfly_C #(.data_width(16)) BF_3_2  (
.A_real( stage3_in_real_2 ),.A_imag( stage3_in_imag_2 ), 
.B_real( stage3_in_real_6 ), .B_imag( stage3_in_imag_6 ),
.W_real(  w8_real  ), .W_imag( w8_imag )
, .clk_MAC(clk_100), .aclr( aclr_s3), .sload(sload_s3) 
,.select( counter_out[1:0]), .O_real(stage3_out_real_2  ), .O_imag( stage3_out_imag_2  ) );  

Butterfly_C #(.data_width(16)) BF_3_3  (
.A_real( stage3_in_real_3 ),.A_imag( stage3_in_imag_3 ), 
.B_real( stage3_in_real_7 ), .B_imag( stage3_in_imag_7 ),
.W_real(  w12_real  ), .W_imag( w12_imag )
, .clk_MAC(clk_100), .aclr( aclr_s3), .sload(sload_s3) 
,.select( counter_out[1:0]), .O_real(stage3_out_real_3  ), .O_imag( stage3_out_imag_3  ) );  

Butterfly_D #(.data_width(16)) BF_3_4  (
.A_real( stage3_in_real_0 ),.A_imag( stage3_in_imag_0 ), 
.B_real( stage3_in_real_4 ), .B_imag( stage3_in_imag_4 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s3), .sload(sload_s3) 
,.select( counter_out[1:0]), .O_real(stage3_out_real_4  ), .O_imag( stage3_out_imag_4  ) );  

Butterfly_D #(.data_width(16)) BF_3_5  (
.A_real( stage3_in_real_1 ),.A_imag( stage3_in_imag_1 ), 
.B_real( stage3_in_real_5 ), .B_imag( stage3_in_imag_5 ),
.W_real(  w4_real  ), .W_imag( w4_imag )
, .clk_MAC(clk_100), .aclr( aclr_s3), .sload(sload_s3) 
,.select( counter_out[1:0]), .O_real(stage3_out_real_5  ), .O_imag( stage3_out_imag_5  ) );  

Butterfly_D #(.data_width(16)) BF_3_6  (
.A_real( stage3_in_real_2 ),.A_imag( stage3_in_imag_2 ), 
.B_real( stage3_in_real_6 ), .B_imag( stage3_in_imag_6 ),
.W_real(  w8_real  ), .W_imag( w8_imag )
, .clk_MAC(clk_100), .aclr( aclr_s3), .sload(sload_s3) 
,.select( counter_out[1:0]), .O_real(stage3_out_real_6  ), .O_imag( stage3_out_imag_6  ) );  

Butterfly_D #(.data_width(16)) BF_3_7  (
.A_real( stage3_in_real_3 ),.A_imag( stage3_in_imag_3 ), 
.B_real( stage3_in_real_7 ), .B_imag( stage3_in_imag_7 ),
.W_real(  w12_real  ), .W_imag( w12_imag )
, .clk_MAC(clk_100), .aclr( aclr_s3), .sload(sload_s3) 
,.select( counter_out[1:0]), .O_real(stage3_out_real_7  ), .O_imag( stage3_out_imag_7  ) );  

/////////////////////////////////////////////////////////////////
Butterfly_C #(.data_width(16)) BF_3_8  (
.A_real( stage3_in_real_8 ),.A_imag( stage3_in_imag_8 ), 
.B_real( stage3_in_real_12 ), .B_imag( stage3_in_imag_12 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s3), .sload(sload_s3) 
,.select( counter_out[1:0]), .O_real(stage3_out_real_8  ), .O_imag( stage3_out_imag_8  ) );  

Butterfly_C #(.data_width(16)) BF_3_9  (
.A_real( stage3_in_real_9 ),.A_imag( stage3_in_imag_9 ), 
.B_real( stage3_in_real_13 ), .B_imag( stage3_in_imag_13 ),
.W_real(  w4_real  ), .W_imag( w4_imag )
, .clk_MAC(clk_100), .aclr( aclr_s3), .sload(sload_s3) 
,.select( counter_out[1:0]), .O_real(stage3_out_real_9  ), .O_imag( stage3_out_imag_9  ) );  

Butterfly_C #(.data_width(16)) BF_3_10  (
.A_real( stage3_in_real_10 ),.A_imag( stage3_in_imag_10 ), 
.B_real( stage3_in_real_14 ), .B_imag( stage3_in_imag_14 ),
.W_real(  w8_real  ), .W_imag( w8_imag )
, .clk_MAC(clk_100), .aclr( aclr_s3), .sload(sload_s3) 
,.select( counter_out[1:0]), .O_real(stage3_out_real_10  ), .O_imag( stage3_out_imag_10  ) );  

Butterfly_C #(.data_width(16)) BF_3_11  (
.A_real( stage3_in_real_11 ),.A_imag( stage3_in_imag_11 ), 
.B_real( stage3_in_real_15 ), .B_imag( stage3_in_imag_15 ),
.W_real(  w12_real  ), .W_imag( w12_imag )
, .clk_MAC(clk_100), .aclr( aclr_s3), .sload(sload_s3) 
,.select( counter_out[1:0]), .O_real(stage3_out_real_11  ), .O_imag( stage3_out_imag_11  ) );  

Butterfly_D #(.data_width(16)) BF_3_12  (
.A_real( stage3_in_real_8 ),.A_imag( stage3_in_imag_8 ), 
.B_real( stage3_in_real_12 ), .B_imag( stage3_in_imag_12 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s3), .sload(sload_s3) 
,.select( counter_out[1:0]), .O_real(stage3_out_real_12  ), .O_imag( stage3_out_imag_12  ) );  

Butterfly_D #(.data_width(16)) BF_3_13  (
.A_real( stage3_in_real_9 ),.A_imag( stage3_in_imag_9 ), 
.B_real( stage3_in_real_13 ), .B_imag( stage3_in_imag_13 ),
.W_real(  w4_real  ), .W_imag( w4_imag )
, .clk_MAC(clk_100), .aclr( aclr_s3), .sload(sload_s3) 
,.select( counter_out[1:0]), .O_real(stage3_out_real_13  ), .O_imag( stage3_out_imag_13  ) );  

Butterfly_D #(.data_width(16)) BF_3_14  (
.A_real( stage3_in_real_10 ),.A_imag( stage3_in_imag_10 ), 
.B_real( stage3_in_real_14 ), .B_imag( stage3_in_imag_14 ),
.W_real(  w8_real  ), .W_imag( w8_imag )
, .clk_MAC(clk_100), .aclr( aclr_s3), .sload(sload_s3) 
,.select( counter_out[1:0]), .O_real(stage3_out_real_14  ), .O_imag( stage3_out_imag_14  ) );  

Butterfly_D #(.data_width(16)) BF_3_15  (
.A_real( stage3_in_real_11 ),.A_imag( stage3_in_imag_11 ), 
.B_real( stage3_in_real_15 ), .B_imag( stage3_in_imag_15 ),
.W_real(  w12_real  ), .W_imag( w12_imag )
, .clk_MAC(clk_100), .aclr( aclr_s3), .sload(sload_s3) 
,.select( counter_out[1:0]), .O_real(stage3_out_real_15  ), .O_imag( stage3_out_imag_15  ) );  

/////////////////////////////////////////////////////////////////
Butterfly_C #(.data_width(16)) BF_3_16  (
.A_real( stage3_in_real_16 ),.A_imag( stage3_in_imag_16 ), 
.B_real( stage3_in_real_20 ), .B_imag( stage3_in_imag_20 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s3), .sload(sload_s3) 
,.select( counter_out[1:0]), .O_real(stage3_out_real_16  ), .O_imag( stage3_out_imag_16  ) );  

Butterfly_C #(.data_width(16)) BF_3_17  (
.A_real( stage3_in_real_17 ),.A_imag( stage3_in_imag_17 ), 
.B_real( stage3_in_real_21 ), .B_imag( stage3_in_imag_21 ),
.W_real(  w4_real  ), .W_imag( w4_imag )
, .clk_MAC(clk_100), .aclr( aclr_s3), .sload(sload_s3) 
,.select( counter_out[1:0]), .O_real(stage3_out_real_17  ), .O_imag( stage3_out_imag_17  ) );  

Butterfly_C #(.data_width(16)) BF_3_18  (
.A_real( stage3_in_real_18 ),.A_imag( stage3_in_imag_18 ), 
.B_real( stage3_in_real_22 ), .B_imag( stage3_in_imag_22 ),
.W_real(  w8_real  ), .W_imag( w8_imag )
, .clk_MAC(clk_100), .aclr( aclr_s3), .sload(sload_s3) 
,.select( counter_out[1:0]), .O_real(stage3_out_real_18  ), .O_imag( stage3_out_imag_18  ) );  

Butterfly_C #(.data_width(16)) BF_3_19  (
.A_real( stage3_in_real_19 ),.A_imag( stage3_in_imag_19 ), 
.B_real( stage3_in_real_23 ), .B_imag( stage3_in_imag_23 ),
.W_real(  w12_real  ), .W_imag( w12_imag )
, .clk_MAC(clk_100), .aclr( aclr_s3), .sload(sload_s3) 
,.select( counter_out[1:0]), .O_real(stage3_out_real_19  ), .O_imag( stage3_out_imag_19  ) );  

Butterfly_D #(.data_width(16)) BF_3_20  (
.A_real( stage3_in_real_16 ),.A_imag( stage3_in_imag_16 ), 
.B_real( stage3_in_real_20 ), .B_imag( stage3_in_imag_20 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s3), .sload(sload_s3) 
,.select( counter_out[1:0]), .O_real(stage3_out_real_20  ), .O_imag( stage3_out_imag_20  ) );  

Butterfly_D #(.data_width(16)) BF_3_21  (
.A_real( stage3_in_real_17 ),.A_imag( stage3_in_imag_17 ), 
.B_real( stage3_in_real_21 ), .B_imag( stage3_in_imag_21 ),
.W_real(  w4_real  ), .W_imag( w4_imag )
, .clk_MAC(clk_100), .aclr( aclr_s3), .sload(sload_s3) 
,.select( counter_out[1:0]), .O_real(stage3_out_real_21  ), .O_imag( stage3_out_imag_21  ) );  

Butterfly_D #(.data_width(16)) BF_3_22  (
.A_real( stage3_in_real_18 ),.A_imag( stage3_in_imag_18 ), 
.B_real( stage3_in_real_22 ), .B_imag( stage3_in_imag_22 ),
.W_real(  w8_real  ), .W_imag( w8_imag )
, .clk_MAC(clk_100), .aclr( aclr_s3), .sload(sload_s3) 
,.select( counter_out[1:0]), .O_real(stage3_out_real_22  ), .O_imag( stage3_out_imag_22  ) );  

Butterfly_D #(.data_width(16)) BF_3_23  (
.A_real( stage3_in_real_19 ),.A_imag( stage3_in_imag_19 ), 
.B_real( stage3_in_real_23 ), .B_imag( stage3_in_imag_23 ),
.W_real(  w12_real  ), .W_imag( w12_imag )
, .clk_MAC(clk_100), .aclr( aclr_s3), .sload(sload_s3) 
,.select( counter_out[1:0]), .O_real(stage3_out_real_23  ), .O_imag( stage3_out_imag_23  ) );  

/////////////////////////////////////////////////////////////////
Butterfly_C #(.data_width(16)) BF_3_24  (
.A_real( stage3_in_real_24 ),.A_imag( stage3_in_imag_24 ), 
.B_real( stage3_in_real_28 ), .B_imag( stage3_in_imag_28 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s3), .sload(sload_s3) 
,.select( counter_out[1:0]), .O_real(stage3_out_real_24  ), .O_imag( stage3_out_imag_24  ) );  

Butterfly_C #(.data_width(16)) BF_3_25  (
.A_real( stage3_in_real_25 ),.A_imag( stage3_in_imag_25 ), 
.B_real( stage3_in_real_29 ), .B_imag( stage3_in_imag_29 ),
.W_real(  w4_real  ), .W_imag( w4_imag )
, .clk_MAC(clk_100), .aclr( aclr_s3), .sload(sload_s3) 
,.select( counter_out[1:0]), .O_real(stage3_out_real_25  ), .O_imag( stage3_out_imag_25  ) );  

Butterfly_C #(.data_width(16)) BF_3_26  (
.A_real( stage3_in_real_26 ),.A_imag( stage3_in_imag_26 ), 
.B_real( stage3_in_real_30 ), .B_imag( stage3_in_imag_30 ),
.W_real(  w8_real  ), .W_imag( w8_imag )
, .clk_MAC(clk_100), .aclr( aclr_s3), .sload(sload_s3) 
,.select( counter_out[1:0]), .O_real(stage3_out_real_26  ), .O_imag( stage3_out_imag_26  ) );  

Butterfly_C #(.data_width(16)) BF_3_27  (
.A_real( stage3_in_real_27 ),.A_imag( stage3_in_imag_27 ), 
.B_real( stage3_in_real_31 ), .B_imag( stage3_in_imag_31 ),
.W_real(  w12_real  ), .W_imag( w12_imag )
, .clk_MAC(clk_100), .aclr( aclr_s3), .sload(sload_s3) 
,.select( counter_out[1:0]), .O_real(stage3_out_real_27  ), .O_imag( stage3_out_imag_27  ) );  

Butterfly_D #(.data_width(16)) BF_3_28  (
.A_real( stage3_in_real_24 ),.A_imag( stage3_in_imag_24 ), 
.B_real( stage3_in_real_28 ), .B_imag( stage3_in_imag_28 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s3), .sload(sload_s3) 
,.select( counter_out[1:0]), .O_real(stage3_out_real_28  ), .O_imag( stage3_out_imag_28  ) );  

Butterfly_D #(.data_width(16)) BF_3_29  (
.A_real( stage3_in_real_25 ),.A_imag( stage3_in_imag_25 ), 
.B_real( stage3_in_real_29 ), .B_imag( stage3_in_imag_29 ),
.W_real(  w4_real  ), .W_imag( w4_imag )
, .clk_MAC(clk_100), .aclr( aclr_s3), .sload(sload_s3) 
,.select( counter_out[1:0]), .O_real(stage3_out_real_29  ), .O_imag( stage3_out_imag_29  ) );  

Butterfly_D #(.data_width(16)) BF_3_30  (
.A_real( stage3_in_real_26 ),.A_imag( stage3_in_imag_26 ), 
.B_real( stage3_in_real_30 ), .B_imag( stage3_in_imag_30 ),
.W_real(  w8_real  ), .W_imag( w8_imag )
, .clk_MAC(clk_100), .aclr( aclr_s3), .sload(sload_s3) 
,.select( counter_out[1:0]), .O_real(stage3_out_real_30  ), .O_imag( stage3_out_imag_30  ) );  

Butterfly_D #(.data_width(16)) BF_3_31  (
.A_real( stage3_in_real_27 ),.A_imag( stage3_in_imag_27 ), 
.B_real( stage3_in_real_31 ), .B_imag( stage3_in_imag_31 ),
.W_real(  w12_real  ), .W_imag( w12_imag )
, .clk_MAC(clk_100), .aclr( aclr_s3), .sload(sload_s3) 
,.select( counter_out[1:0]), .O_real(stage3_out_real_31  ), .O_imag( stage3_out_imag_31  ) );  

/////////////////////////////////////////////////////////////////


Butterfly_C #(.data_width(16)) BF_4_0  (
.A_real( stage4_in_real_0 ),.A_imag(stage4_in_imag_0), 
.B_real( stage4_in_real_8 ), .B_imag(  stage4_in_imag_8 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s4), .sload(sload_s4) 
,.select( counter_out[1:0]), .O_real(stage4_out_real_0  ), .O_imag( stage4_out_imag_0  ) );  

Butterfly_C #(.data_width(16)) BF_4_1  (
.A_real( stage4_in_real_1 ),.A_imag(stage4_in_imag_1), 
.B_real( stage4_in_real_9 ), .B_imag(  stage4_in_imag_9 ),
.W_real(  w2_real  ), .W_imag( w2_imag )
, .clk_MAC(clk_100), .aclr( aclr_s4), .sload(sload_s4) 
,.select( counter_out[1:0]), .O_real(stage4_out_real_1  ), .O_imag( stage4_out_imag_1  ) );  

Butterfly_C #(.data_width(16)) BF_4_2  (
.A_real( stage4_in_real_2 ),.A_imag(stage4_in_imag_2), 
.B_real( stage4_in_real_10 ), .B_imag(  stage4_in_imag_10 ),
.W_real(  w4_real  ), .W_imag( w4_imag )
, .clk_MAC(clk_100), .aclr( aclr_s4), .sload(sload_s4) 
,.select( counter_out[1:0]), .O_real(stage4_out_real_2  ), .O_imag( stage4_out_imag_2  ) );  

Butterfly_C #(.data_width(16)) BF_4_3  (
.A_real( stage4_in_real_3 ),.A_imag(stage4_in_imag_3), 
.B_real( stage4_in_real_11 ), .B_imag(  stage4_in_imag_11 ),
.W_real(  w6_real  ), .W_imag( w6_imag )
, .clk_MAC(clk_100), .aclr( aclr_s4), .sload(sload_s4) 
,.select( counter_out[1:0]), .O_real(stage4_out_real_3  ), .O_imag( stage4_out_imag_3  ) );  

Butterfly_C #(.data_width(16)) BF_4_4  (
.A_real( stage4_in_real_4 ),.A_imag(stage4_in_imag_4), 
.B_real( stage4_in_real_12 ), .B_imag(  stage4_in_imag_12 ),
.W_real(  w8_real  ), .W_imag( w8_imag )
, .clk_MAC(clk_100), .aclr( aclr_s4), .sload(sload_s4) 
,.select( counter_out[1:0]), .O_real(stage4_out_real_4  ), .O_imag( stage4_out_imag_4  ) );  

Butterfly_C #(.data_width(16)) BF_4_5  (
.A_real( stage4_in_real_5 ),.A_imag(stage4_in_imag_5), 
.B_real( stage4_in_real_13 ), .B_imag(  stage4_in_imag_13 ),
.W_real(  w14_real  ), .W_imag( w10_imag )
, .clk_MAC(clk_100), .aclr( aclr_s4), .sload(sload_s4) 
,.select( counter_out[1:0]), .O_real(stage4_out_real_5  ), .O_imag( stage4_out_imag_5  ) );  

Butterfly_C #(.data_width(16)) BF_4_6  (
.A_real( stage4_in_real_6 ),.A_imag(stage4_in_imag_6), 
.B_real( stage4_in_real_14 ), .B_imag(  stage4_in_imag_14 ),
.W_real(  w12_real  ), .W_imag( w12_imag )
, .clk_MAC(clk_100), .aclr( aclr_s4), .sload(sload_s4) 
,.select( counter_out[1:0]), .O_real(stage4_out_real_6  ), .O_imag( stage4_out_imag_6  ) );  

Butterfly_C #(.data_width(16)) BF_4_7  (
.A_real( stage4_in_real_7 ),.A_imag(stage4_in_imag_7), 
.B_real( stage4_in_real_15 ), .B_imag(  stage4_in_imag_15 ),
.W_real(  w14_real  ), .W_imag( w14_imag )
, .clk_MAC(clk_100), .aclr( aclr_s4), .sload(sload_s4) 
,.select( counter_out[1:0]), .O_real(stage4_out_real_7  ), .O_imag( stage4_out_imag_7  ) );  

Butterfly_D #(.data_width(16)) BF_4_8  (
.A_real( stage4_in_real_0 ),.A_imag(stage4_in_imag_0), 
.B_real( stage4_in_real_8 ), .B_imag(  stage4_in_imag_8 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s4), .sload(sload_s4) 
,.select( counter_out[1:0]), .O_real(stage4_out_real_8  ), .O_imag( stage4_out_imag_8  ) );  

Butterfly_D #(.data_width(16)) BF_4_9  (
.A_real( stage4_in_real_1 ),.A_imag(stage4_in_imag_1), 
.B_real( stage4_in_real_9 ), .B_imag(  stage4_in_imag_9 ),
.W_real(  w2_real  ), .W_imag( w2_imag )
, .clk_MAC(clk_100), .aclr( aclr_s4), .sload(sload_s4) 
,.select( counter_out[1:0]), .O_real(stage4_out_real_9  ), .O_imag( stage4_out_imag_9  ) );  

Butterfly_D #(.data_width(16)) BF_4_10  (
.A_real( stage4_in_real_2 ),.A_imag(stage4_in_imag_2), 
.B_real( stage4_in_real_10 ), .B_imag(  stage4_in_imag_10 ),
.W_real(  w4_real  ), .W_imag( w4_imag )
, .clk_MAC(clk_100), .aclr( aclr_s4), .sload(sload_s4) 
,.select( counter_out[1:0]), .O_real(stage4_out_real_10  ), .O_imag( stage4_out_imag_10  ) );  

Butterfly_D #(.data_width(16)) BF_4_11  (
.A_real( stage4_in_real_3 ),.A_imag(stage4_in_imag_3), 
.B_real( stage4_in_real_11 ), .B_imag(  stage4_in_imag_11 ),
.W_real(  w6_real  ), .W_imag( w6_imag )
, .clk_MAC(clk_100), .aclr( aclr_s4), .sload(sload_s4) 
,.select( counter_out[1:0]), .O_real(stage4_out_real_11  ), .O_imag( stage4_out_imag_11  ) );  

Butterfly_D #(.data_width(16)) BF_4_12  (
.A_real( stage4_in_real_4 ),.A_imag(stage4_in_imag_4), 
.B_real( stage4_in_real_12 ), .B_imag(  stage4_in_imag_12 ),
.W_real(  w8_real  ), .W_imag( w8_imag )
, .clk_MAC(clk_100), .aclr( aclr_s4), .sload(sload_s4) 
,.select( counter_out[1:0]), .O_real(stage4_out_real_12  ), .O_imag( stage4_out_imag_12  ) );  

Butterfly_D #(.data_width(16)) BF_4_13  (
.A_real( stage4_in_real_5 ),.A_imag(stage4_in_imag_5), 
.B_real( stage4_in_real_13 ), .B_imag(  stage4_in_imag_13 ),
.W_real( w14_real  ), .W_imag( w10_imag )
, .clk_MAC(clk_100), .aclr( aclr_s4), .sload(sload_s4) 
,.select( counter_out[1:0]), .O_real(stage4_out_real_13  ), .O_imag( stage4_out_imag_13  ) );  

Butterfly_D #(.data_width(16)) BF_4_14  (
.A_real( stage4_in_real_6 ),.A_imag(stage4_in_imag_6), 
.B_real( stage4_in_real_14 ), .B_imag(  stage4_in_imag_14 ),
.W_real(  w12_real  ), .W_imag( w12_imag )
, .clk_MAC(clk_100), .aclr( aclr_s4), .sload(sload_s4) 
,.select( counter_out[1:0]), .O_real(stage4_out_real_14  ), .O_imag( stage4_out_imag_14  ) );  

Butterfly_D #(.data_width(16)) BF_4_15  (
.A_real( stage4_in_real_7 ),.A_imag(stage4_in_imag_7), 
.B_real( stage4_in_real_15 ), .B_imag(  stage4_in_imag_15 ),
.W_real(  w14_real  ), .W_imag( w14_imag )
, .clk_MAC(clk_100), .aclr( aclr_s4), .sload(sload_s4) 
,.select( counter_out[1:0]), .O_real(stage4_out_real_15  ), .O_imag( stage4_out_imag_15  ) );  

/////////////////////////////////////////////////////////////////
Butterfly_C #(.data_width(16)) BF_4_16  (
.A_real( stage4_in_real_16 ),.A_imag(stage4_in_imag_16), 
.B_real( stage4_in_real_24 ), .B_imag(  stage4_in_imag_24 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s4), .sload(sload_s4) 
,.select( counter_out[1:0]), .O_real(stage4_out_real_16  ), .O_imag( stage4_out_imag_16  ) );  

Butterfly_C #(.data_width(16)) BF_4_17  (
.A_real( stage4_in_real_17 ),.A_imag(stage4_in_imag_17), 
.B_real( stage4_in_real_25 ), .B_imag(  stage4_in_imag_25 ),
.W_real(  w2_real  ), .W_imag( w2_imag )
, .clk_MAC(clk_100), .aclr( aclr_s4), .sload(sload_s4) 
,.select( counter_out[1:0]), .O_real(stage4_out_real_17  ), .O_imag( stage4_out_imag_17  ) );  

Butterfly_C #(.data_width(16)) BF_4_18  (
.A_real( stage4_in_real_18 ),.A_imag(stage4_in_imag_18), 
.B_real( stage4_in_real_26 ), .B_imag(  stage4_in_imag_26 ),
.W_real(  w4_real  ), .W_imag( w4_imag )
, .clk_MAC(clk_100), .aclr( aclr_s4), .sload(sload_s4) 
,.select( counter_out[1:0]), .O_real(stage4_out_real_18  ), .O_imag( stage4_out_imag_18  ) );  

Butterfly_C #(.data_width(16)) BF_4_19  (
.A_real( stage4_in_real_19 ),.A_imag(stage4_in_imag_19), 
.B_real( stage4_in_real_27 ), .B_imag(  stage4_in_imag_27 ),
.W_real(  w6_real  ), .W_imag( w6_imag )
, .clk_MAC(clk_100), .aclr( aclr_s4), .sload(sload_s4) 
,.select( counter_out[1:0]), .O_real(stage4_out_real_19  ), .O_imag( stage4_out_imag_19  ) );  

Butterfly_C #(.data_width(16)) BF_4_20  (
.A_real( stage4_in_real_20 ),.A_imag(stage4_in_imag_20), 
.B_real( stage4_in_real_28 ), .B_imag(  stage4_in_imag_28 ),
.W_real(  w8_real  ), .W_imag( w8_imag )
, .clk_MAC(clk_100), .aclr( aclr_s4), .sload(sload_s4) 
,.select( counter_out[1:0]), .O_real(stage4_out_real_20  ), .O_imag( stage4_out_imag_20  ) );  

Butterfly_C #(.data_width(16)) BF_4_21  (
.A_real( stage4_in_real_21 ),.A_imag(stage4_in_imag_21), 
.B_real( stage4_in_real_29 ), .B_imag(  stage4_in_imag_29 ),
.W_real(  w14_real  ), .W_imag( w10_imag )
, .clk_MAC(clk_100), .aclr( aclr_s4), .sload(sload_s4) 
,.select( counter_out[1:0]), .O_real(stage4_out_real_21  ), .O_imag( stage4_out_imag_21  ) );  

Butterfly_C #(.data_width(16)) BF_4_22  (
.A_real( stage4_in_real_22 ),.A_imag(stage4_in_imag_22), 
.B_real( stage4_in_real_30 ), .B_imag(  stage4_in_imag_30 ),
.W_real(  w12_real  ), .W_imag( w12_imag )
, .clk_MAC(clk_100), .aclr( aclr_s4), .sload(sload_s4) 
,.select( counter_out[1:0]), .O_real(stage4_out_real_22  ), .O_imag( stage4_out_imag_22  ) );  

Butterfly_C #(.data_width(16)) BF_4_23  (
.A_real( stage4_in_real_23 ),.A_imag(stage4_in_imag_23), 
.B_real( stage4_in_real_31 ), .B_imag(  stage4_in_imag_31 ),
.W_real(  w14_real  ), .W_imag( w14_imag )
, .clk_MAC(clk_100), .aclr( aclr_s4), .sload(sload_s4) 
,.select( counter_out[1:0]), .O_real(stage4_out_real_23  ), .O_imag( stage4_out_imag_23  ) );  

Butterfly_D #(.data_width(16)) BF_4_24  (
.A_real( stage4_in_real_16 ),.A_imag(stage4_in_imag_16), 
.B_real( stage4_in_real_24 ), .B_imag(  stage4_in_imag_24 ),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s4), .sload(sload_s4) 
,.select( counter_out[1:0]), .O_real(stage4_out_real_24  ), .O_imag( stage4_out_imag_24  ) );  

Butterfly_D #(.data_width(16)) BF_4_25  (
.A_real( stage4_in_real_17 ),.A_imag(stage4_in_imag_17), 
.B_real( stage4_in_real_25 ), .B_imag(  stage4_in_imag_25 ),
.W_real(  w2_real  ), .W_imag( w2_imag )
, .clk_MAC(clk_100), .aclr( aclr_s4), .sload(sload_s4) 
,.select( counter_out[1:0]), .O_real(stage4_out_real_25  ), .O_imag( stage4_out_imag_25  ) );  

Butterfly_D #(.data_width(16)) BF_4_26  (
.A_real( stage4_in_real_18 ),.A_imag(stage4_in_imag_18), 
.B_real( stage4_in_real_26 ), .B_imag(  stage4_in_imag_26 ),
.W_real(  w4_real  ), .W_imag( w4_imag )
, .clk_MAC(clk_100), .aclr( aclr_s4), .sload(sload_s4) 
,.select( counter_out[1:0]), .O_real(stage4_out_real_26  ), .O_imag( stage4_out_imag_26  ) );  

Butterfly_D #(.data_width(16)) BF_4_27  (
.A_real( stage4_in_real_19 ),.A_imag(stage4_in_imag_19), 
.B_real( stage4_in_real_27 ), .B_imag(  stage4_in_imag_27 ),
.W_real(  w6_real  ), .W_imag( w6_imag )
, .clk_MAC(clk_100), .aclr( aclr_s4), .sload(sload_s4) 
,.select( counter_out[1:0]), .O_real(stage4_out_real_27  ), .O_imag( stage4_out_imag_27  ) );  

Butterfly_D #(.data_width(16)) BF_4_28  (
.A_real( stage4_in_real_20 ),.A_imag(stage4_in_imag_20), 
.B_real( stage4_in_real_28 ), .B_imag(  stage4_in_imag_28 ),
.W_real(  w8_real  ), .W_imag( w8_imag )
, .clk_MAC(clk_100), .aclr( aclr_s4), .sload(sload_s4) 
,.select( counter_out[1:0]), .O_real(stage4_out_real_28  ), .O_imag( stage4_out_imag_28  ) );  

Butterfly_D #(.data_width(16)) BF_4_29  (
.A_real( stage4_in_real_21 ),.A_imag(stage4_in_imag_21), 
.B_real( stage4_in_real_29 ), .B_imag(  stage4_in_imag_29 ),
.W_real( w14_real  ), .W_imag( w10_imag )
, .clk_MAC(clk_100), .aclr( aclr_s4), .sload(sload_s4) 
,.select( counter_out[1:0]), .O_real(stage4_out_real_29  ), .O_imag( stage4_out_imag_29  ) );  

Butterfly_D #(.data_width(16)) BF_4_30  (
.A_real( stage4_in_real_22 ),.A_imag(stage4_in_imag_22), 
.B_real( stage4_in_real_30 ), .B_imag(  stage4_in_imag_30 ),
.W_real(  w12_real  ), .W_imag( w12_imag )
, .clk_MAC(clk_100), .aclr( aclr_s4), .sload(sload_s4) 
,.select( counter_out[1:0]), .O_real(stage4_out_real_30  ), .O_imag( stage4_out_imag_30  ) );  

Butterfly_D #(.data_width(16)) BF_4_31  (
.A_real( stage4_in_real_23 ),.A_imag(stage4_in_imag_23), 
.B_real( stage4_in_real_31 ), .B_imag(  stage4_in_imag_31 ),
.W_real(  w14_real  ), .W_imag( w14_imag )
, .clk_MAC(clk_100), .aclr( aclr_s4), .sload(sload_s4) 
,.select( counter_out[1:0]), .O_real(stage4_out_real_31  ), .O_imag( stage4_out_imag_31  ) );  

/////////////////////////////////////////////////////////////////



Butterfly_C #(.data_width(16)) BF_5_0  (
.A_real( stage5_in_real_0),.A_imag(stage5_in_imag_0), 
.B_real( stage5_in_real_16), .B_imag(  stage5_in_imag_16),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s5), .sload(sload_s5) 
,.select( counter_out[1:0]), .O_real(stage5_out_real_0  ), .O_imag( stage5_out_imag_0  ) );  

Butterfly_C #(.data_width(16)) BF_5_1  (
.A_real( stage5_in_real_1),.A_imag(stage5_in_imag_1), 
.B_real( stage5_in_real_17), .B_imag(  stage5_in_imag_17),
.W_real(  w1_real  ), .W_imag( w1_imag )
, .clk_MAC(clk_100), .aclr( aclr_s5), .sload(sload_s5) 
,.select( counter_out[1:0]), .O_real(stage5_out_real_1  ), .O_imag( stage5_out_imag_1  ) );  

Butterfly_C #(.data_width(16)) BF_5_2  (
.A_real( stage5_in_real_2),.A_imag(stage5_in_imag_2), 
.B_real( stage5_in_real_18), .B_imag(  stage5_in_imag_18),
.W_real(  w2_real  ), .W_imag( w2_imag )
, .clk_MAC(clk_100), .aclr( aclr_s5), .sload(sload_s5) 
,.select( counter_out[1:0]), .O_real(stage5_out_real_2  ), .O_imag( stage5_out_imag_2  ) );  

Butterfly_C #(.data_width(16)) BF_5_3  (
.A_real( stage5_in_real_3),.A_imag(stage5_in_imag_3), 
.B_real( stage5_in_real_19), .B_imag(  stage5_in_imag_19),
.W_real(  w3_real  ), .W_imag( w3_imag )
, .clk_MAC(clk_100), .aclr( aclr_s5), .sload(sload_s5) 
,.select( counter_out[1:0]), .O_real(stage5_out_real_3  ), .O_imag( stage5_out_imag_3  ) );  

Butterfly_C #(.data_width(16)) BF_5_4  (
.A_real( stage5_in_real_4),.A_imag(stage5_in_imag_4), 
.B_real( stage5_in_real_20), .B_imag(  stage5_in_imag_20),
.W_real(  w4_real  ), .W_imag( w4_imag )
, .clk_MAC(clk_100), .aclr( aclr_s5), .sload(sload_s5) 
,.select( counter_out[1:0]), .O_real(stage5_out_real_4  ), .O_imag( stage5_out_imag_4  ) );  

Butterfly_C #(.data_width(16)) BF_5_5  (
.A_real( stage5_in_real_5),.A_imag(stage5_in_imag_5), 
.B_real( stage5_in_real_21), .B_imag(  stage5_in_imag_21),
.W_real(  w5_real  ), .W_imag( w5_imag )
, .clk_MAC(clk_100), .aclr( aclr_s5), .sload(sload_s5) 
,.select( counter_out[1:0]), .O_real(stage5_out_real_5  ), .O_imag( stage5_out_imag_5  ) );  

Butterfly_C #(.data_width(16)) BF_5_6  (
.A_real( stage5_in_real_6),.A_imag(stage5_in_imag_6), 
.B_real( stage5_in_real_22), .B_imag(  stage5_in_imag_22),
.W_real(  w6_real  ), .W_imag( w6_imag )
, .clk_MAC(clk_100), .aclr( aclr_s5), .sload(sload_s5) 
,.select( counter_out[1:0]), .O_real(stage5_out_real_6  ), .O_imag( stage5_out_imag_6  ) );  

Butterfly_C #(.data_width(16)) BF_5_7  (
.A_real( stage5_in_real_7),.A_imag(stage5_in_imag_7), 
.B_real( stage5_in_real_23), .B_imag(  stage5_in_imag_23),
.W_real(  w7_real  ), .W_imag( w7_imag )
, .clk_MAC(clk_100), .aclr( aclr_s5), .sload(sload_s5) 
,.select( counter_out[1:0]), .O_real(stage5_out_real_7  ), .O_imag( stage5_out_imag_7  ) );  

Butterfly_C #(.data_width(16)) BF_5_8  (
.A_real( stage5_in_real_8),.A_imag(stage5_in_imag_8), 
.B_real( stage5_in_real_24), .B_imag(  stage5_in_imag_24),
.W_real(  w8_real  ), .W_imag( w8_imag )
, .clk_MAC(clk_100), .aclr( aclr_s5), .sload(sload_s5) 
,.select( counter_out[1:0]), .O_real(stage5_out_real_8  ), .O_imag( stage5_out_imag_8  ) );  

Butterfly_C #(.data_width(16)) BF_5_9  (
.A_real( stage5_in_real_9),.A_imag(stage5_in_imag_9), 
.B_real( stage5_in_real_25), .B_imag(  stage5_in_imag_25),
.W_real(  w9_real  ), .W_imag( w9_imag )
, .clk_MAC(clk_100), .aclr( aclr_s5), .sload(sload_s5) 
,.select( counter_out[1:0]), .O_real(stage5_out_real_9  ), .O_imag( stage5_out_imag_9  ) );  

Butterfly_C #(.data_width(16)) BF_5_10  (
.A_real( stage5_in_real_10),.A_imag(stage5_in_imag_10), 
.B_real( stage5_in_real_26), .B_imag(  stage5_in_imag_26),
.W_real(  w10_real  ), .W_imag( w10_imag )
, .clk_MAC(clk_100), .aclr( aclr_s5), .sload(sload_s5) 
,.select( counter_out[1:0]), .O_real(stage5_out_real_10  ), .O_imag( stage5_out_imag_10  ) );  

Butterfly_C #(.data_width(16)) BF_5_11  (
.A_real( stage5_in_real_11),.A_imag(stage5_in_imag_11), 
.B_real( stage5_in_real_27), .B_imag(  stage5_in_imag_27),
.W_real(  w11_real  ), .W_imag( w11_imag )
, .clk_MAC(clk_100), .aclr( aclr_s5), .sload(sload_s5) 
,.select( counter_out[1:0]), .O_real(stage5_out_real_11  ), .O_imag( stage5_out_imag_11  ) );  

Butterfly_C #(.data_width(16)) BF_5_12  (
.A_real( stage5_in_real_12),.A_imag(stage5_in_imag_12), 
.B_real( stage5_in_real_28), .B_imag(  stage5_in_imag_28),
.W_real(  w12_real  ), .W_imag( w12_imag )
, .clk_MAC(clk_100), .aclr( aclr_s5), .sload(sload_s5) 
,.select( counter_out[1:0]), .O_real(stage5_out_real_12  ), .O_imag( stage5_out_imag_12  ) );  

Butterfly_C #(.data_width(16)) BF_5_13  (
.A_real( stage5_in_real_13),.A_imag(stage5_in_imag_13), 
.B_real( stage5_in_real_29), .B_imag(  stage5_in_imag_29),
.W_real( w13_real  ), .W_imag( w13_imag )
, .clk_MAC(clk_100), .aclr( aclr_s5), .sload(sload_s5) 
,.select( counter_out[1:0]), .O_real(stage5_out_real_13  ), .O_imag( stage5_out_imag_13  ) );  

Butterfly_C #(.data_width(16)) BF_5_14  (
.A_real( stage5_in_real_14),.A_imag(stage5_in_imag_14), 
.B_real( stage5_in_real_30), .B_imag(  stage5_in_imag_30),
.W_real(  w14_real  ), .W_imag( w14_imag )
, .clk_MAC(clk_100), .aclr( aclr_s5), .sload(sload_s5) 
,.select( counter_out[1:0]), .O_real(stage5_out_real_14  ), .O_imag( stage5_out_imag_14  ) );  

Butterfly_C #(.data_width(16)) BF_5_15  (
.A_real( stage5_in_real_15),.A_imag(stage5_in_imag_15), 
.B_real( stage5_in_real_31), .B_imag(  stage5_in_imag_31),
.W_real(  w15_real  ), .W_imag( w15_imag )
, .clk_MAC(clk_100), .aclr( aclr_s5), .sload(sload_s5) 
,.select( counter_out[1:0]), .O_real(stage5_out_real_15  ), .O_imag( stage5_out_imag_15  ) );  

Butterfly_D #(.data_width(16)) BF_5_16  (
.A_real( stage5_in_real_0),.A_imag(stage5_in_imag_0), 
.B_real( stage5_in_real_16), .B_imag(  stage5_in_imag_16),
.W_real(  w0_real  ), .W_imag( w0_imag )
, .clk_MAC(clk_100), .aclr( aclr_s5), .sload(sload_s5) 
,.select( counter_out[1:0]), .O_real(stage5_out_real_16  ), .O_imag( stage5_out_imag_16  ) );  

Butterfly_D #(.data_width(16)) BF_5_17  (
.A_real( stage5_in_real_1),.A_imag(stage5_in_imag_1), 
.B_real( stage5_in_real_17), .B_imag(  stage5_in_imag_17),
.W_real(  w1_real  ), .W_imag( w1_imag )
, .clk_MAC(clk_100), .aclr( aclr_s5), .sload(sload_s5) 
,.select( counter_out[1:0]), .O_real(stage5_out_real_17  ), .O_imag( stage5_out_imag_17  ) );  

Butterfly_D #(.data_width(16)) BF_5_18  (
.A_real( stage5_in_real_2),.A_imag(stage5_in_imag_2), 
.B_real( stage5_in_real_18), .B_imag(  stage5_in_imag_18),
.W_real(  w2_real  ), .W_imag( w2_imag )
, .clk_MAC(clk_100), .aclr( aclr_s5), .sload(sload_s5) 
,.select( counter_out[1:0]), .O_real(stage5_out_real_18  ), .O_imag( stage5_out_imag_18  ) );  

Butterfly_D #(.data_width(16)) BF_5_19  (
.A_real( stage5_in_real_3),.A_imag(stage5_in_imag_3), 
.B_real( stage5_in_real_19), .B_imag(  stage5_in_imag_19),
.W_real(  w3_real  ), .W_imag( w3_imag )
, .clk_MAC(clk_100), .aclr( aclr_s5), .sload(sload_s5) 
,.select( counter_out[1:0]), .O_real(stage5_out_real_19  ), .O_imag( stage5_out_imag_19  ) );  

Butterfly_D #(.data_width(16)) BF_5_20  (
.A_real( stage5_in_real_4),.A_imag(stage5_in_imag_4), 
.B_real( stage5_in_real_20), .B_imag(  stage5_in_imag_20),
.W_real(  w4_real  ), .W_imag( w4_imag )
, .clk_MAC(clk_100), .aclr( aclr_s5), .sload(sload_s5) 
,.select( counter_out[1:0]), .O_real(stage5_out_real_20  ), .O_imag( stage5_out_imag_20  ) );  

Butterfly_D #(.data_width(16)) BF_5_21  (
.A_real( stage5_in_real_5),.A_imag(stage5_in_imag_5), 
.B_real( stage5_in_real_21), .B_imag(  stage5_in_imag_21),
.W_real(  w5_real  ), .W_imag( w5_imag )
, .clk_MAC(clk_100), .aclr( aclr_s5), .sload(sload_s5) 
,.select( counter_out[1:0]), .O_real(stage5_out_real_21  ), .O_imag( stage5_out_imag_21  ) );  

Butterfly_D #(.data_width(16)) BF_5_22  (
.A_real( stage5_in_real_6),.A_imag(stage5_in_imag_6), 
.B_real( stage5_in_real_22), .B_imag(  stage5_in_imag_22),
.W_real( w6_real  ), .W_imag( w6_imag )
, .clk_MAC(clk_100), .aclr( aclr_s5), .sload(sload_s5) 
,.select( counter_out[1:0]), .O_real(stage5_out_real_22  ), .O_imag( stage5_out_imag_22  ) );  

Butterfly_D #(.data_width(16)) BF_5_23  (
.A_real( stage5_in_real_7),.A_imag(stage5_in_imag_7), 
.B_real( stage5_in_real_23), .B_imag(  stage5_in_imag_23),
.W_real(  w7_real  ), .W_imag( w7_imag )
, .clk_MAC(clk_100), .aclr( aclr_s5), .sload(sload_s5) 
,.select( counter_out[1:0]), .O_real(stage5_out_real_23  ), .O_imag( stage5_out_imag_23  ) );  

Butterfly_D #(.data_width(16)) BF_5_24  (
.A_real( stage5_in_real_8),.A_imag(stage5_in_imag_8), 
.B_real( stage5_in_real_24), .B_imag(  stage5_in_imag_24),
.W_real(  w8_real  ), .W_imag( w8_imag )
, .clk_MAC(clk_100), .aclr( aclr_s5), .sload(sload_s5) 
,.select( counter_out[1:0]), .O_real(stage5_out_real_24  ), .O_imag( stage5_out_imag_24  ) );  

Butterfly_D #(.data_width(16)) BF_5_25  (
.A_real( stage5_in_real_9),.A_imag(stage5_in_imag_9), 
.B_real( stage5_in_real_25), .B_imag(  stage5_in_imag_25),
.W_real( w9_real  ), .W_imag( w9_imag )
, .clk_MAC(clk_100), .aclr( aclr_s5), .sload(sload_s5) 
,.select( counter_out[1:0]), .O_real(stage5_out_real_25  ), .O_imag( stage5_out_imag_25  ) );  

Butterfly_D #(.data_width(16)) BF_5_26  (
.A_real( stage5_in_real_10),.A_imag(stage5_in_imag_10), 
.B_real( stage5_in_real_26), .B_imag(  stage5_in_imag_26),
.W_real(  w10_real  ), .W_imag( w10_imag )
, .clk_MAC(clk_100), .aclr( aclr_s5), .sload(sload_s5) 
,.select( counter_out[1:0]), .O_real(stage5_out_real_26  ), .O_imag( stage5_out_imag_26  ) );  

Butterfly_D #(.data_width(16)) BF_5_27  (
.A_real( stage5_in_real_11),.A_imag(stage5_in_imag_11), 
.B_real( stage5_in_real_27), .B_imag(  stage5_in_imag_27),
.W_real(  w11_real  ), .W_imag( w11_imag )
, .clk_MAC(clk_100), .aclr( aclr_s5), .sload(sload_s5) 
,.select( counter_out[1:0]), .O_real(stage5_out_real_27  ), .O_imag( stage5_out_imag_27  ) );  

Butterfly_D #(.data_width(16)) BF_5_28  (
.A_real( stage5_in_real_12),.A_imag(stage5_in_imag_12), 
.B_real( stage5_in_real_28), .B_imag(  stage5_in_imag_28),
.W_real(  w12_real  ), .W_imag( w12_imag )
, .clk_MAC(clk_100), .aclr( aclr_s5), .sload(sload_s5) 
,.select( counter_out[1:0]), .O_real(stage5_out_real_28  ), .O_imag( stage5_out_imag_28  ) );  

Butterfly_D #(.data_width(16)) BF_5_29  (
.A_real( stage5_in_real_13),.A_imag(stage5_in_imag_13), 
.B_real( stage5_in_real_29), .B_imag(  stage5_in_imag_29),
.W_real( w13_real  ), .W_imag( w13_imag )
, .clk_MAC(clk_100), .aclr( aclr_s5), .sload(sload_s5) 
,.select( counter_out[1:0]), .O_real(stage5_out_real_29  ), .O_imag( stage5_out_imag_29  ) );  

Butterfly_D #(.data_width(16)) BF_5_30  (
.A_real( stage5_in_real_14),.A_imag(stage5_in_imag_14), 
.B_real( stage5_in_real_30), .B_imag(  stage5_in_imag_30),
.W_real( w14_real  ), .W_imag( w14_imag )
, .clk_MAC(clk_100), .aclr( aclr_s5), .sload(sload_s5) 
,.select( counter_out[1:0]), .O_real(stage5_out_real_30  ), .O_imag( stage5_out_imag_30  ) );  

Butterfly_D #(.data_width(16)) BF_5_31  (
.A_real( stage5_in_real_15),.A_imag(stage5_in_imag_15), 
.B_real( stage5_in_real_31), .B_imag(  stage5_in_imag_31),
.W_real(  w15_real  ), .W_imag( w15_imag )
, .clk_MAC(clk_100), .aclr( aclr_s5), .sload(sload_s5) 
,.select( counter_out[1:0]), .O_real(stage5_out_real_31  ), .O_imag( stage5_out_imag_31  ) );  

//////////////////////////////////////////////////////////////////////////////////////////////////////////////////////

/////////////////////////////////////////////////////////////////

reg signed [15:0] stage1_in_r_real_0;
reg signed [15:0] stage1_in_r_imag_0;
reg signed [15:0] stage1_in_r_real_1;
reg signed [15:0] stage1_in_r_imag_1;
reg signed [15:0] stage1_in_r_real_2;
reg signed [15:0] stage1_in_r_imag_2;
reg signed [15:0] stage1_in_r_real_3;
reg signed [15:0] stage1_in_r_imag_3;
reg signed [15:0] stage1_in_r_real_4;
reg signed [15:0] stage1_in_r_imag_4;
reg signed [15:0] stage1_in_r_real_5;
reg signed [15:0] stage1_in_r_imag_5;
reg signed [15:0] stage1_in_r_real_6;
reg signed [15:0] stage1_in_r_imag_6;
reg signed [15:0] stage1_in_r_real_7;
reg signed [15:0] stage1_in_r_imag_7;
reg signed [15:0] stage1_in_r_real_8;
reg signed [15:0] stage1_in_r_imag_8;
reg signed [15:0] stage1_in_r_real_9;
reg signed [15:0] stage1_in_r_imag_9;
reg signed [15:0] stage1_in_r_real_10;
reg signed [15:0] stage1_in_r_imag_10;
reg signed [15:0] stage1_in_r_real_11;
reg signed [15:0] stage1_in_r_imag_11;
reg signed [15:0] stage1_in_r_real_12;
reg signed [15:0] stage1_in_r_imag_12;
reg signed [15:0] stage1_in_r_real_13;
reg signed [15:0] stage1_in_r_imag_13;
reg signed [15:0] stage1_in_r_real_14;
reg signed [15:0] stage1_in_r_imag_14;
reg signed [15:0] stage1_in_r_real_15;
reg signed [15:0] stage1_in_r_imag_15;
reg signed [15:0] stage1_in_r_real_16;
reg signed [15:0] stage1_in_r_imag_16;
reg signed [15:0] stage1_in_r_real_17;
reg signed [15:0] stage1_in_r_imag_17;
reg signed [15:0] stage1_in_r_real_18;
reg signed [15:0] stage1_in_r_imag_18;
reg signed [15:0] stage1_in_r_real_19;
reg signed [15:0] stage1_in_r_imag_19;
reg signed [15:0] stage1_in_r_real_20;
reg signed [15:0] stage1_in_r_imag_20;
reg signed [15:0] stage1_in_r_real_21;
reg signed [15:0] stage1_in_r_imag_21;
reg signed [15:0] stage1_in_r_real_22;
reg signed [15:0] stage1_in_r_imag_22;
reg signed [15:0] stage1_in_r_real_23;
reg signed [15:0] stage1_in_r_imag_23;
reg signed [15:0] stage1_in_r_real_24;
reg signed [15:0] stage1_in_r_imag_24;
reg signed [15:0] stage1_in_r_real_25;
reg signed [15:0] stage1_in_r_imag_25;
reg signed [15:0] stage1_in_r_real_26;
reg signed [15:0] stage1_in_r_imag_26;
reg signed [15:0] stage1_in_r_real_27;
reg signed [15:0] stage1_in_r_imag_27;
reg signed [15:0] stage1_in_r_real_28;
reg signed [15:0] stage1_in_r_imag_28;
reg signed [15:0] stage1_in_r_real_29;
reg signed [15:0] stage1_in_r_imag_29;
reg signed [15:0] stage1_in_r_real_30;
reg signed [15:0] stage1_in_r_imag_30;
reg signed [15:0] stage1_in_r_real_31;
reg signed [15:0] stage1_in_r_imag_31;
reg signed [15:0] stage2_in_r_real_0;
reg signed [15:0] stage2_in_r_imag_0;
reg signed [15:0] stage2_in_r_real_1;
reg signed [15:0] stage2_in_r_imag_1;
reg signed [15:0] stage2_in_r_real_2;
reg signed [15:0] stage2_in_r_imag_2;
reg signed [15:0] stage2_in_r_real_3;
reg signed [15:0] stage2_in_r_imag_3;
reg signed [15:0] stage2_in_r_real_4;
reg signed [15:0] stage2_in_r_imag_4;
reg signed [15:0] stage2_in_r_real_5;
reg signed [15:0] stage2_in_r_imag_5;
reg signed [15:0] stage2_in_r_real_6;
reg signed [15:0] stage2_in_r_imag_6;
reg signed [15:0] stage2_in_r_real_7;
reg signed [15:0] stage2_in_r_imag_7;
reg signed [15:0] stage2_in_r_real_8;
reg signed [15:0] stage2_in_r_imag_8;
reg signed [15:0] stage2_in_r_real_9;
reg signed [15:0] stage2_in_r_imag_9;
reg signed [15:0] stage2_in_r_real_10;
reg signed [15:0] stage2_in_r_imag_10;
reg signed [15:0] stage2_in_r_real_11;
reg signed [15:0] stage2_in_r_imag_11;
reg signed [15:0] stage2_in_r_real_12;
reg signed [15:0] stage2_in_r_imag_12;
reg signed [15:0] stage2_in_r_real_13;
reg signed [15:0] stage2_in_r_imag_13;
reg signed [15:0] stage2_in_r_real_14;
reg signed [15:0] stage2_in_r_imag_14;
reg signed [15:0] stage2_in_r_real_15;
reg signed [15:0] stage2_in_r_imag_15;
reg signed [15:0] stage2_in_r_real_16;
reg signed [15:0] stage2_in_r_imag_16;
reg signed [15:0] stage2_in_r_real_17;
reg signed [15:0] stage2_in_r_imag_17;
reg signed [15:0] stage2_in_r_real_18;
reg signed [15:0] stage2_in_r_imag_18;
reg signed [15:0] stage2_in_r_real_19;
reg signed [15:0] stage2_in_r_imag_19;
reg signed [15:0] stage2_in_r_real_20;
reg signed [15:0] stage2_in_r_imag_20;
reg signed [15:0] stage2_in_r_real_21;
reg signed [15:0] stage2_in_r_imag_21;
reg signed [15:0] stage2_in_r_real_22;
reg signed [15:0] stage2_in_r_imag_22;
reg signed [15:0] stage2_in_r_real_23;
reg signed [15:0] stage2_in_r_imag_23;
reg signed [15:0] stage2_in_r_real_24;
reg signed [15:0] stage2_in_r_imag_24;
reg signed [15:0] stage2_in_r_real_25;
reg signed [15:0] stage2_in_r_imag_25;
reg signed [15:0] stage2_in_r_real_26;
reg signed [15:0] stage2_in_r_imag_26;
reg signed [15:0] stage2_in_r_real_27;
reg signed [15:0] stage2_in_r_imag_27;
reg signed [15:0] stage2_in_r_real_28;
reg signed [15:0] stage2_in_r_imag_28;
reg signed [15:0] stage2_in_r_real_29;
reg signed [15:0] stage2_in_r_imag_29;
reg signed [15:0] stage2_in_r_real_30;
reg signed [15:0] stage2_in_r_imag_30;
reg signed [15:0] stage2_in_r_real_31;
reg signed [15:0] stage2_in_r_imag_31;
reg signed [15:0] stage3_in_r_real_0;
reg signed [15:0] stage3_in_r_imag_0;
reg signed [15:0] stage3_in_r_real_1;
reg signed [15:0] stage3_in_r_imag_1;
reg signed [15:0] stage3_in_r_real_2;
reg signed [15:0] stage3_in_r_imag_2;
reg signed [15:0] stage3_in_r_real_3;
reg signed [15:0] stage3_in_r_imag_3;
reg signed [15:0] stage3_in_r_real_4;
reg signed [15:0] stage3_in_r_imag_4;
reg signed [15:0] stage3_in_r_real_5;
reg signed [15:0] stage3_in_r_imag_5;
reg signed [15:0] stage3_in_r_real_6;
reg signed [15:0] stage3_in_r_imag_6;
reg signed [15:0] stage3_in_r_real_7;
reg signed [15:0] stage3_in_r_imag_7;
reg signed [15:0] stage3_in_r_real_8;
reg signed [15:0] stage3_in_r_imag_8;
reg signed [15:0] stage3_in_r_real_9;
reg signed [15:0] stage3_in_r_imag_9;
reg signed [15:0] stage3_in_r_real_10;
reg signed [15:0] stage3_in_r_imag_10;
reg signed [15:0] stage3_in_r_real_11;
reg signed [15:0] stage3_in_r_imag_11;
reg signed [15:0] stage3_in_r_real_12;
reg signed [15:0] stage3_in_r_imag_12;
reg signed [15:0] stage3_in_r_real_13;
reg signed [15:0] stage3_in_r_imag_13;
reg signed [15:0] stage3_in_r_real_14;
reg signed [15:0] stage3_in_r_imag_14;
reg signed [15:0] stage3_in_r_real_15;
reg signed [15:0] stage3_in_r_imag_15;
reg signed [15:0] stage3_in_r_real_16;
reg signed [15:0] stage3_in_r_imag_16;
reg signed [15:0] stage3_in_r_real_17;
reg signed [15:0] stage3_in_r_imag_17;
reg signed [15:0] stage3_in_r_real_18;
reg signed [15:0] stage3_in_r_imag_18;
reg signed [15:0] stage3_in_r_real_19;
reg signed [15:0] stage3_in_r_imag_19;
reg signed [15:0] stage3_in_r_real_20;
reg signed [15:0] stage3_in_r_imag_20;
reg signed [15:0] stage3_in_r_real_21;
reg signed [15:0] stage3_in_r_imag_21;
reg signed [15:0] stage3_in_r_real_22;
reg signed [15:0] stage3_in_r_imag_22;
reg signed [15:0] stage3_in_r_real_23;
reg signed [15:0] stage3_in_r_imag_23;
reg signed [15:0] stage3_in_r_real_24;
reg signed [15:0] stage3_in_r_imag_24;
reg signed [15:0] stage3_in_r_real_25;
reg signed [15:0] stage3_in_r_imag_25;
reg signed [15:0] stage3_in_r_real_26;
reg signed [15:0] stage3_in_r_imag_26;
reg signed [15:0] stage3_in_r_real_27;
reg signed [15:0] stage3_in_r_imag_27;
reg signed [15:0] stage3_in_r_real_28;
reg signed [15:0] stage3_in_r_imag_28;
reg signed [15:0] stage3_in_r_real_29;
reg signed [15:0] stage3_in_r_imag_29;
reg signed [15:0] stage3_in_r_real_30;
reg signed [15:0] stage3_in_r_imag_30;
reg signed [15:0] stage3_in_r_real_31;
reg signed [15:0] stage3_in_r_imag_31;
reg signed [15:0] stage4_in_r_real_0;
reg signed [15:0] stage4_in_r_imag_0;
reg signed [15:0] stage4_in_r_real_1;
reg signed [15:0] stage4_in_r_imag_1;
reg signed [15:0] stage4_in_r_real_2;
reg signed [15:0] stage4_in_r_imag_2;
reg signed [15:0] stage4_in_r_real_3;
reg signed [15:0] stage4_in_r_imag_3;
reg signed [15:0] stage4_in_r_real_4;
reg signed [15:0] stage4_in_r_imag_4;
reg signed [15:0] stage4_in_r_real_5;
reg signed [15:0] stage4_in_r_imag_5;
reg signed [15:0] stage4_in_r_real_6;
reg signed [15:0] stage4_in_r_imag_6;
reg signed [15:0] stage4_in_r_real_7;
reg signed [15:0] stage4_in_r_imag_7;
reg signed [15:0] stage4_in_r_real_8;
reg signed [15:0] stage4_in_r_imag_8;
reg signed [15:0] stage4_in_r_real_9;
reg signed [15:0] stage4_in_r_imag_9;
reg signed [15:0] stage4_in_r_real_10;
reg signed [15:0] stage4_in_r_imag_10;
reg signed [15:0] stage4_in_r_real_11;
reg signed [15:0] stage4_in_r_imag_11;
reg signed [15:0] stage4_in_r_real_12;
reg signed [15:0] stage4_in_r_imag_12;
reg signed [15:0] stage4_in_r_real_13;
reg signed [15:0] stage4_in_r_imag_13;
reg signed [15:0] stage4_in_r_real_14;
reg signed [15:0] stage4_in_r_imag_14;
reg signed [15:0] stage4_in_r_real_15;
reg signed [15:0] stage4_in_r_imag_15;
reg signed [15:0] stage4_in_r_real_16;
reg signed [15:0] stage4_in_r_imag_16;
reg signed [15:0] stage4_in_r_real_17;
reg signed [15:0] stage4_in_r_imag_17;
reg signed [15:0] stage4_in_r_real_18;
reg signed [15:0] stage4_in_r_imag_18;
reg signed [15:0] stage4_in_r_real_19;
reg signed [15:0] stage4_in_r_imag_19;
reg signed [15:0] stage4_in_r_real_20;
reg signed [15:0] stage4_in_r_imag_20;
reg signed [15:0] stage4_in_r_real_21;
reg signed [15:0] stage4_in_r_imag_21;
reg signed [15:0] stage4_in_r_real_22;
reg signed [15:0] stage4_in_r_imag_22;
reg signed [15:0] stage4_in_r_real_23;
reg signed [15:0] stage4_in_r_imag_23;
reg signed [15:0] stage4_in_r_real_24;
reg signed [15:0] stage4_in_r_imag_24;
reg signed [15:0] stage4_in_r_real_25;
reg signed [15:0] stage4_in_r_imag_25;
reg signed [15:0] stage4_in_r_real_26;
reg signed [15:0] stage4_in_r_imag_26;
reg signed [15:0] stage4_in_r_real_27;
reg signed [15:0] stage4_in_r_imag_27;
reg signed [15:0] stage4_in_r_real_28;
reg signed [15:0] stage4_in_r_imag_28;
reg signed [15:0] stage4_in_r_real_29;
reg signed [15:0] stage4_in_r_imag_29;
reg signed [15:0] stage4_in_r_real_30;
reg signed [15:0] stage4_in_r_imag_30;
reg signed [15:0] stage4_in_r_real_31;
reg signed [15:0] stage4_in_r_imag_31;
reg signed [15:0] stage5_in_r_real_0;
reg signed [15:0] stage5_in_r_imag_0;
reg signed [15:0] stage5_in_r_real_1;
reg signed [15:0] stage5_in_r_imag_1;
reg signed [15:0] stage5_in_r_real_2;
reg signed [15:0] stage5_in_r_imag_2;
reg signed [15:0] stage5_in_r_real_3;
reg signed [15:0] stage5_in_r_imag_3;
reg signed [15:0] stage5_in_r_real_4;
reg signed [15:0] stage5_in_r_imag_4;
reg signed [15:0] stage5_in_r_real_5;
reg signed [15:0] stage5_in_r_imag_5;
reg signed [15:0] stage5_in_r_real_6;
reg signed [15:0] stage5_in_r_imag_6;
reg signed [15:0] stage5_in_r_real_7;
reg signed [15:0] stage5_in_r_imag_7;
reg signed [15:0] stage5_in_r_real_8;
reg signed [15:0] stage5_in_r_imag_8;
reg signed [15:0] stage5_in_r_real_9;
reg signed [15:0] stage5_in_r_imag_9;
reg signed [15:0] stage5_in_r_real_10;
reg signed [15:0] stage5_in_r_imag_10;
reg signed [15:0] stage5_in_r_real_11;
reg signed [15:0] stage5_in_r_imag_11;
reg signed [15:0] stage5_in_r_real_12;
reg signed [15:0] stage5_in_r_imag_12;
reg signed [15:0] stage5_in_r_real_13;
reg signed [15:0] stage5_in_r_imag_13;
reg signed [15:0] stage5_in_r_real_14;
reg signed [15:0] stage5_in_r_imag_14;
reg signed [15:0] stage5_in_r_real_15;
reg signed [15:0] stage5_in_r_imag_15;
reg signed [15:0] stage5_in_r_real_16;
reg signed [15:0] stage5_in_r_imag_16;
reg signed [15:0] stage5_in_r_real_17;
reg signed [15:0] stage5_in_r_imag_17;
reg signed [15:0] stage5_in_r_real_18;
reg signed [15:0] stage5_in_r_imag_18;
reg signed [15:0] stage5_in_r_real_19;
reg signed [15:0] stage5_in_r_imag_19;
reg signed [15:0] stage5_in_r_real_20;
reg signed [15:0] stage5_in_r_imag_20;
reg signed [15:0] stage5_in_r_real_21;
reg signed [15:0] stage5_in_r_imag_21;
reg signed [15:0] stage5_in_r_real_22;
reg signed [15:0] stage5_in_r_imag_22;
reg signed [15:0] stage5_in_r_real_23;
reg signed [15:0] stage5_in_r_imag_23;
reg signed [15:0] stage5_in_r_real_24;
reg signed [15:0] stage5_in_r_imag_24;
reg signed [15:0] stage5_in_r_real_25;
reg signed [15:0] stage5_in_r_imag_25;
reg signed [15:0] stage5_in_r_real_26;
reg signed [15:0] stage5_in_r_imag_26;
reg signed [15:0] stage5_in_r_real_27;
reg signed [15:0] stage5_in_r_imag_27;
reg signed [15:0] stage5_in_r_real_28;
reg signed [15:0] stage5_in_r_imag_28;
reg signed [15:0] stage5_in_r_real_29;
reg signed [15:0] stage5_in_r_imag_29;
reg signed [15:0] stage5_in_r_real_30;
reg signed [15:0] stage5_in_r_imag_30;
reg signed [15:0] stage5_in_r_real_31;
reg signed [15:0] stage5_in_r_imag_31;

//[31:0] >> all stages except stage5
assign stage1_in_real_0  = stage1_in_r_real_0;
assign stage1_in_imag_0  = stage1_in_r_imag_0;
assign stage1_in_real_1  = stage1_in_r_real_1;
assign stage1_in_imag_1  = stage1_in_r_imag_1;
assign stage1_in_real_2  = stage1_in_r_real_2;
assign stage1_in_imag_2  = stage1_in_r_imag_2;
assign stage1_in_real_3  = stage1_in_r_real_3;
assign stage1_in_imag_3  = stage1_in_r_imag_3;
assign stage1_in_real_4  = stage1_in_r_real_4;
assign stage1_in_imag_4  = stage1_in_r_imag_4;
assign stage1_in_real_5  = stage1_in_r_real_5;
assign stage1_in_imag_5  = stage1_in_r_imag_5;
assign stage1_in_real_6  = stage1_in_r_real_6;
assign stage1_in_imag_6  = stage1_in_r_imag_6;
assign stage1_in_real_7  = stage1_in_r_real_7;
assign stage1_in_imag_7  = stage1_in_r_imag_7;
assign stage1_in_real_8  = stage1_in_r_real_8;
assign stage1_in_imag_8  = stage1_in_r_imag_8;
assign stage1_in_real_9  = stage1_in_r_real_9;
assign stage1_in_imag_9  = stage1_in_r_imag_9;
assign stage1_in_real_10  = stage1_in_r_real_10;
assign stage1_in_imag_10  = stage1_in_r_imag_10;
assign stage1_in_real_11  = stage1_in_r_real_11;
assign stage1_in_imag_11  = stage1_in_r_imag_11;
assign stage1_in_real_12  = stage1_in_r_real_12;
assign stage1_in_imag_12  = stage1_in_r_imag_12;
assign stage1_in_real_13  = stage1_in_r_real_13;
assign stage1_in_imag_13  = stage1_in_r_imag_13;
assign stage1_in_real_14  = stage1_in_r_real_14;
assign stage1_in_imag_14  = stage1_in_r_imag_14;
assign stage1_in_real_15  = stage1_in_r_real_15;
assign stage1_in_imag_15  = stage1_in_r_imag_15;
assign stage1_in_real_16  = stage1_in_r_real_16;
assign stage1_in_imag_16  = stage1_in_r_imag_16;
assign stage1_in_real_17  = stage1_in_r_real_17;
assign stage1_in_imag_17  = stage1_in_r_imag_17;
assign stage1_in_real_18  = stage1_in_r_real_18;
assign stage1_in_imag_18  = stage1_in_r_imag_18;
assign stage1_in_real_19  = stage1_in_r_real_19;
assign stage1_in_imag_19  = stage1_in_r_imag_19;
assign stage1_in_real_20  = stage1_in_r_real_20;
assign stage1_in_imag_20  = stage1_in_r_imag_20;
assign stage1_in_real_21  = stage1_in_r_real_21;
assign stage1_in_imag_21  = stage1_in_r_imag_21;
assign stage1_in_real_22  = stage1_in_r_real_22;
assign stage1_in_imag_22  = stage1_in_r_imag_22;
assign stage1_in_real_23  = stage1_in_r_real_23;
assign stage1_in_imag_23  = stage1_in_r_imag_23;
assign stage1_in_real_24  = stage1_in_r_real_24;
assign stage1_in_imag_24  = stage1_in_r_imag_24;
assign stage1_in_real_25  = stage1_in_r_real_25;
assign stage1_in_imag_25  = stage1_in_r_imag_25;
assign stage1_in_real_26  = stage1_in_r_real_26;
assign stage1_in_imag_26  = stage1_in_r_imag_26;
assign stage1_in_real_27  = stage1_in_r_real_27;
assign stage1_in_imag_27  = stage1_in_r_imag_27;
assign stage1_in_real_28  = stage1_in_r_real_28;
assign stage1_in_imag_28  = stage1_in_r_imag_28;
assign stage1_in_real_29  = stage1_in_r_real_29;
assign stage1_in_imag_29  = stage1_in_r_imag_29;
assign stage1_in_real_30  = stage1_in_r_real_30;
assign stage1_in_imag_30  = stage1_in_r_imag_30;
assign stage1_in_real_31  = stage1_in_r_real_31;
assign stage1_in_imag_31  = stage1_in_r_imag_31;
assign stage2_in_real_0  = stage2_in_r_real_0;
assign stage2_in_imag_0  = stage2_in_r_imag_0;
assign stage2_in_real_1  = stage2_in_r_real_1;
assign stage2_in_imag_1  = stage2_in_r_imag_1;
assign stage2_in_real_2  = stage2_in_r_real_2;
assign stage2_in_imag_2  = stage2_in_r_imag_2;
assign stage2_in_real_3  = stage2_in_r_real_3;
assign stage2_in_imag_3  = stage2_in_r_imag_3;
assign stage2_in_real_4  = stage2_in_r_real_4;
assign stage2_in_imag_4  = stage2_in_r_imag_4;
assign stage2_in_real_5  = stage2_in_r_real_5;
assign stage2_in_imag_5  = stage2_in_r_imag_5;
assign stage2_in_real_6  = stage2_in_r_real_6;
assign stage2_in_imag_6  = stage2_in_r_imag_6;
assign stage2_in_real_7  = stage2_in_r_real_7;
assign stage2_in_imag_7  = stage2_in_r_imag_7;
assign stage2_in_real_8  = stage2_in_r_real_8;
assign stage2_in_imag_8  = stage2_in_r_imag_8;
assign stage2_in_real_9  = stage2_in_r_real_9;
assign stage2_in_imag_9  = stage2_in_r_imag_9;
assign stage2_in_real_10  = stage2_in_r_real_10;
assign stage2_in_imag_10  = stage2_in_r_imag_10;
assign stage2_in_real_11  = stage2_in_r_real_11;
assign stage2_in_imag_11  = stage2_in_r_imag_11;
assign stage2_in_real_12  = stage2_in_r_real_12;
assign stage2_in_imag_12  = stage2_in_r_imag_12;
assign stage2_in_real_13  = stage2_in_r_real_13;
assign stage2_in_imag_13  = stage2_in_r_imag_13;
assign stage2_in_real_14  = stage2_in_r_real_14;
assign stage2_in_imag_14  = stage2_in_r_imag_14;
assign stage2_in_real_15  = stage2_in_r_real_15;
assign stage2_in_imag_15  = stage2_in_r_imag_15;
assign stage2_in_real_16  = stage2_in_r_real_16;
assign stage2_in_imag_16  = stage2_in_r_imag_16;
assign stage2_in_real_17  = stage2_in_r_real_17;
assign stage2_in_imag_17  = stage2_in_r_imag_17;
assign stage2_in_real_18  = stage2_in_r_real_18;
assign stage2_in_imag_18  = stage2_in_r_imag_18;
assign stage2_in_real_19  = stage2_in_r_real_19;
assign stage2_in_imag_19  = stage2_in_r_imag_19;
assign stage2_in_real_20  = stage2_in_r_real_20;
assign stage2_in_imag_20  = stage2_in_r_imag_20;
assign stage2_in_real_21  = stage2_in_r_real_21;
assign stage2_in_imag_21  = stage2_in_r_imag_21;
assign stage2_in_real_22  = stage2_in_r_real_22;
assign stage2_in_imag_22  = stage2_in_r_imag_22;
assign stage2_in_real_23  = stage2_in_r_real_23;
assign stage2_in_imag_23  = stage2_in_r_imag_23;
assign stage2_in_real_24  = stage2_in_r_real_24;
assign stage2_in_imag_24  = stage2_in_r_imag_24;
assign stage2_in_real_25  = stage2_in_r_real_25;
assign stage2_in_imag_25  = stage2_in_r_imag_25;
assign stage2_in_real_26  = stage2_in_r_real_26;
assign stage2_in_imag_26  = stage2_in_r_imag_26;
assign stage2_in_real_27  = stage2_in_r_real_27;
assign stage2_in_imag_27  = stage2_in_r_imag_27;
assign stage2_in_real_28  = stage2_in_r_real_28;
assign stage2_in_imag_28  = stage2_in_r_imag_28;
assign stage2_in_real_29  = stage2_in_r_real_29;
assign stage2_in_imag_29  = stage2_in_r_imag_29;
assign stage2_in_real_30  = stage2_in_r_real_30;
assign stage2_in_imag_30  = stage2_in_r_imag_30;
assign stage2_in_real_31  = stage2_in_r_real_31;
assign stage2_in_imag_31  = stage2_in_r_imag_31;
assign stage3_in_real_0  = stage3_in_r_real_0;
assign stage3_in_imag_0  = stage3_in_r_imag_0;
assign stage3_in_real_1  = stage3_in_r_real_1;
assign stage3_in_imag_1  = stage3_in_r_imag_1;
assign stage3_in_real_2  = stage3_in_r_real_2;
assign stage3_in_imag_2  = stage3_in_r_imag_2;
assign stage3_in_real_3  = stage3_in_r_real_3;
assign stage3_in_imag_3  = stage3_in_r_imag_3;
assign stage3_in_real_4  = stage3_in_r_real_4;
assign stage3_in_imag_4  = stage3_in_r_imag_4;
assign stage3_in_real_5  = stage3_in_r_real_5;
assign stage3_in_imag_5  = stage3_in_r_imag_5;
assign stage3_in_real_6  = stage3_in_r_real_6;
assign stage3_in_imag_6  = stage3_in_r_imag_6;
assign stage3_in_real_7  = stage3_in_r_real_7;
assign stage3_in_imag_7  = stage3_in_r_imag_7;
assign stage3_in_real_8  = stage3_in_r_real_8;
assign stage3_in_imag_8  = stage3_in_r_imag_8;
assign stage3_in_real_9  = stage3_in_r_real_9;
assign stage3_in_imag_9  = stage3_in_r_imag_9;
assign stage3_in_real_10  = stage3_in_r_real_10;
assign stage3_in_imag_10  = stage3_in_r_imag_10;
assign stage3_in_real_11  = stage3_in_r_real_11;
assign stage3_in_imag_11  = stage3_in_r_imag_11;
assign stage3_in_real_12  = stage3_in_r_real_12;
assign stage3_in_imag_12  = stage3_in_r_imag_12;
assign stage3_in_real_13  = stage3_in_r_real_13;
assign stage3_in_imag_13  = stage3_in_r_imag_13;
assign stage3_in_real_14  = stage3_in_r_real_14;
assign stage3_in_imag_14  = stage3_in_r_imag_14;
assign stage3_in_real_15  = stage3_in_r_real_15;
assign stage3_in_imag_15  = stage3_in_r_imag_15;
assign stage3_in_real_16  = stage3_in_r_real_16;
assign stage3_in_imag_16  = stage3_in_r_imag_16;
assign stage3_in_real_17  = stage3_in_r_real_17;
assign stage3_in_imag_17  = stage3_in_r_imag_17;
assign stage3_in_real_18  = stage3_in_r_real_18;
assign stage3_in_imag_18  = stage3_in_r_imag_18;
assign stage3_in_real_19  = stage3_in_r_real_19;
assign stage3_in_imag_19  = stage3_in_r_imag_19;
assign stage3_in_real_20  = stage3_in_r_real_20;
assign stage3_in_imag_20  = stage3_in_r_imag_20;
assign stage3_in_real_21  = stage3_in_r_real_21;
assign stage3_in_imag_21  = stage3_in_r_imag_21;
assign stage3_in_real_22  = stage3_in_r_real_22;
assign stage3_in_imag_22  = stage3_in_r_imag_22;
assign stage3_in_real_23  = stage3_in_r_real_23;
assign stage3_in_imag_23  = stage3_in_r_imag_23;
assign stage3_in_real_24  = stage3_in_r_real_24;
assign stage3_in_imag_24  = stage3_in_r_imag_24;
assign stage3_in_real_25  = stage3_in_r_real_25;
assign stage3_in_imag_25  = stage3_in_r_imag_25;
assign stage3_in_real_26  = stage3_in_r_real_26;
assign stage3_in_imag_26  = stage3_in_r_imag_26;
assign stage3_in_real_27  = stage3_in_r_real_27;
assign stage3_in_imag_27  = stage3_in_r_imag_27;
assign stage3_in_real_28  = stage3_in_r_real_28;
assign stage3_in_imag_28  = stage3_in_r_imag_28;
assign stage3_in_real_29  = stage3_in_r_real_29;
assign stage3_in_imag_29  = stage3_in_r_imag_29;
assign stage3_in_real_30  = stage3_in_r_real_30;
assign stage3_in_imag_30  = stage3_in_r_imag_30;
assign stage3_in_real_31  = stage3_in_r_real_31;
assign stage3_in_imag_31  = stage3_in_r_imag_31;
assign stage4_in_real_0  = stage4_in_r_real_0;
assign stage4_in_imag_0  = stage4_in_r_imag_0;
assign stage4_in_real_1  = stage4_in_r_real_1;
assign stage4_in_imag_1  = stage4_in_r_imag_1;
assign stage4_in_real_2  = stage4_in_r_real_2;
assign stage4_in_imag_2  = stage4_in_r_imag_2;
assign stage4_in_real_3  = stage4_in_r_real_3;
assign stage4_in_imag_3  = stage4_in_r_imag_3;
assign stage4_in_real_4  = stage4_in_r_real_4;
assign stage4_in_imag_4  = stage4_in_r_imag_4;
assign stage4_in_real_5  = stage4_in_r_real_5;
assign stage4_in_imag_5  = stage4_in_r_imag_5;
assign stage4_in_real_6  = stage4_in_r_real_6;
assign stage4_in_imag_6  = stage4_in_r_imag_6;
assign stage4_in_real_7  = stage4_in_r_real_7;
assign stage4_in_imag_7  = stage4_in_r_imag_7;
assign stage4_in_real_8  = stage4_in_r_real_8;
assign stage4_in_imag_8  = stage4_in_r_imag_8;
assign stage4_in_real_9  = stage4_in_r_real_9;
assign stage4_in_imag_9  = stage4_in_r_imag_9;
assign stage4_in_real_10  = stage4_in_r_real_10;
assign stage4_in_imag_10  = stage4_in_r_imag_10;
assign stage4_in_real_11  = stage4_in_r_real_11;
assign stage4_in_imag_11  = stage4_in_r_imag_11;
assign stage4_in_real_12  = stage4_in_r_real_12;
assign stage4_in_imag_12  = stage4_in_r_imag_12;
assign stage4_in_real_13  = stage4_in_r_real_13;
assign stage4_in_imag_13  = stage4_in_r_imag_13;
assign stage4_in_real_14  = stage4_in_r_real_14;
assign stage4_in_imag_14  = stage4_in_r_imag_14;
assign stage4_in_real_15  = stage4_in_r_real_15;
assign stage4_in_imag_15  = stage4_in_r_imag_15;
assign stage4_in_real_16  = stage4_in_r_real_16;
assign stage4_in_imag_16  = stage4_in_r_imag_16;
assign stage4_in_real_17  = stage4_in_r_real_17;
assign stage4_in_imag_17  = stage4_in_r_imag_17;
assign stage4_in_real_18  = stage4_in_r_real_18;
assign stage4_in_imag_18  = stage4_in_r_imag_18;
assign stage4_in_real_19  = stage4_in_r_real_19;
assign stage4_in_imag_19  = stage4_in_r_imag_19;
assign stage4_in_real_20  = stage4_in_r_real_20;
assign stage4_in_imag_20  = stage4_in_r_imag_20;
assign stage4_in_real_21  = stage4_in_r_real_21;
assign stage4_in_imag_21  = stage4_in_r_imag_21;
assign stage4_in_real_22  = stage4_in_r_real_22;
assign stage4_in_imag_22  = stage4_in_r_imag_22;
assign stage4_in_real_23  = stage4_in_r_real_23;
assign stage4_in_imag_23  = stage4_in_r_imag_23;
assign stage4_in_real_24  = stage4_in_r_real_24;
assign stage4_in_imag_24  = stage4_in_r_imag_24;
assign stage4_in_real_25  = stage4_in_r_real_25;
assign stage4_in_imag_25  = stage4_in_r_imag_25;
assign stage4_in_real_26  = stage4_in_r_real_26;
assign stage4_in_imag_26  = stage4_in_r_imag_26;
assign stage4_in_real_27  = stage4_in_r_real_27;
assign stage4_in_imag_27  = stage4_in_r_imag_27;
assign stage4_in_real_28  = stage4_in_r_real_28;
assign stage4_in_imag_28  = stage4_in_r_imag_28;
assign stage4_in_real_29  = stage4_in_r_real_29;
assign stage4_in_imag_29  = stage4_in_r_imag_29;
assign stage4_in_real_30  = stage4_in_r_real_30;
assign stage4_in_imag_30  = stage4_in_r_imag_30;
assign stage4_in_real_31  = stage4_in_r_real_31;
assign stage4_in_imag_31  = stage4_in_r_imag_31;



assign stage5_in_real_0  = stage5_in_r_real_0;
assign stage5_in_imag_0  = stage5_in_r_imag_0;
assign stage5_in_real_1  = stage5_in_r_real_1;
assign stage5_in_imag_1  = stage5_in_r_imag_1;
assign stage5_in_real_2  = stage5_in_r_real_2;
assign stage5_in_imag_2  = stage5_in_r_imag_2;
assign stage5_in_real_3  = stage5_in_r_real_3;
assign stage5_in_imag_3  = stage5_in_r_imag_3;
assign stage5_in_real_4  = stage5_in_r_real_4;
assign stage5_in_imag_4  = stage5_in_r_imag_4;
assign stage5_in_real_5  = stage5_in_r_real_5;
assign stage5_in_imag_5  = stage5_in_r_imag_5;
assign stage5_in_real_6  = stage5_in_r_real_6;
assign stage5_in_imag_6  = stage5_in_r_imag_6;
assign stage5_in_real_7  = stage5_in_r_real_7;
assign stage5_in_imag_7  = stage5_in_r_imag_7;
assign stage5_in_real_8  = stage5_in_r_real_8;
assign stage5_in_imag_8  = stage5_in_r_imag_8;
assign stage5_in_real_9  = stage5_in_r_real_9;
assign stage5_in_imag_9  = stage5_in_r_imag_9;
assign stage5_in_real_10  = stage5_in_r_real_10;
assign stage5_in_imag_10  = stage5_in_r_imag_10;
assign stage5_in_real_11  = stage5_in_r_real_11;
assign stage5_in_imag_11  = stage5_in_r_imag_11;
assign stage5_in_real_12  = stage5_in_r_real_12;
assign stage5_in_imag_12  = stage5_in_r_imag_12;
assign stage5_in_real_13  = stage5_in_r_real_13;
assign stage5_in_imag_13  = stage5_in_r_imag_13;
assign stage5_in_real_14  = stage5_in_r_real_14;
assign stage5_in_imag_14  = stage5_in_r_imag_14;
assign stage5_in_real_15  = stage5_in_r_real_15;
assign stage5_in_imag_15  = stage5_in_r_imag_15;
assign stage5_in_real_16  = stage5_in_r_real_16;
assign stage5_in_imag_16  = stage5_in_r_imag_16;
assign stage5_in_real_17  = stage5_in_r_real_17;
assign stage5_in_imag_17  = stage5_in_r_imag_17;
assign stage5_in_real_18  = stage5_in_r_real_18;
assign stage5_in_imag_18  = stage5_in_r_imag_18;
assign stage5_in_real_19  = stage5_in_r_real_19;
assign stage5_in_imag_19  = stage5_in_r_imag_19;
assign stage5_in_real_20  = stage5_in_r_real_20;
assign stage5_in_imag_20  = stage5_in_r_imag_20;
assign stage5_in_real_21  = stage5_in_r_real_21;
assign stage5_in_imag_21  = stage5_in_r_imag_21;
assign stage5_in_real_22  = stage5_in_r_real_22;
assign stage5_in_imag_22  = stage5_in_r_imag_22;
assign stage5_in_real_23  = stage5_in_r_real_23;
assign stage5_in_imag_23  = stage5_in_r_imag_23;
assign stage5_in_real_24  = stage5_in_r_real_24;
assign stage5_in_imag_24  = stage5_in_r_imag_24;
assign stage5_in_real_25  = stage5_in_r_real_25;
assign stage5_in_imag_25  = stage5_in_r_imag_25;
assign stage5_in_real_26  = stage5_in_r_real_26;
assign stage5_in_imag_26  = stage5_in_r_imag_26;
assign stage5_in_real_27  = stage5_in_r_real_27;
assign stage5_in_imag_27  = stage5_in_r_imag_27;
assign stage5_in_real_28  = stage5_in_r_real_28;
assign stage5_in_imag_28  = stage5_in_r_imag_28;
assign stage5_in_real_29  = stage5_in_r_real_29;
assign stage5_in_imag_29  = stage5_in_r_imag_29;
assign stage5_in_real_30  = stage5_in_r_real_30;
assign stage5_in_imag_30  = stage5_in_r_imag_30;
assign stage5_in_real_31  = stage5_in_r_real_31;
assign stage5_in_imag_31  = stage5_in_r_imag_31;


 always @ (posedge clk_20) begin


stage2_in_r_real_0 <= stage1_out_real_0;
stage2_in_r_imag_0  <= stage1_out_imag_0;
stage2_in_r_real_1 <= stage1_out_real_1;
stage2_in_r_imag_1  <= stage1_out_imag_1;
stage2_in_r_real_2 <= stage1_out_real_2;
stage2_in_r_imag_2  <= stage1_out_imag_2;
stage2_in_r_real_3 <= stage1_out_real_3;
stage2_in_r_imag_3  <= stage1_out_imag_3;
stage2_in_r_real_4 <= stage1_out_real_4;
stage2_in_r_imag_4  <= stage1_out_imag_4;
stage2_in_r_real_5 <= stage1_out_real_5;
stage2_in_r_imag_5  <= stage1_out_imag_5;
stage2_in_r_real_6 <= stage1_out_real_6;
stage2_in_r_imag_6  <= stage1_out_imag_6;
stage2_in_r_real_7 <= stage1_out_real_7;
stage2_in_r_imag_7  <= stage1_out_imag_7;
stage2_in_r_real_8 <= stage1_out_real_8;
stage2_in_r_imag_8  <= stage1_out_imag_8;
stage2_in_r_real_9 <= stage1_out_real_9;
stage2_in_r_imag_9  <= stage1_out_imag_9;
stage2_in_r_real_10 <= stage1_out_real_10;
stage2_in_r_imag_10  <= stage1_out_imag_10;
stage2_in_r_real_11 <= stage1_out_real_11;
stage2_in_r_imag_11  <= stage1_out_imag_11;
stage2_in_r_real_12 <= stage1_out_real_12;
stage2_in_r_imag_12  <= stage1_out_imag_12;
stage2_in_r_real_13 <= stage1_out_real_13;
stage2_in_r_imag_13  <= stage1_out_imag_13;
stage2_in_r_real_14 <= stage1_out_real_14;
stage2_in_r_imag_14  <= stage1_out_imag_14;
stage2_in_r_real_15 <= stage1_out_real_15;
stage2_in_r_imag_15  <= stage1_out_imag_15;
stage2_in_r_real_16 <= stage1_out_real_16;
stage2_in_r_imag_16  <= stage1_out_imag_16;
stage2_in_r_real_17 <= stage1_out_real_17;
stage2_in_r_imag_17  <= stage1_out_imag_17;
stage2_in_r_real_18 <= stage1_out_real_18;
stage2_in_r_imag_18  <= stage1_out_imag_18;
stage2_in_r_real_19 <= stage1_out_real_19;
stage2_in_r_imag_19  <= stage1_out_imag_19;
stage2_in_r_real_20 <= stage1_out_real_20;
stage2_in_r_imag_20  <= stage1_out_imag_20;
stage2_in_r_real_21 <= stage1_out_real_21;
stage2_in_r_imag_21  <= stage1_out_imag_21;
stage2_in_r_real_22 <= stage1_out_real_22;
stage2_in_r_imag_22  <= stage1_out_imag_22;
stage2_in_r_real_23 <= stage1_out_real_23;
stage2_in_r_imag_23  <= stage1_out_imag_23;
stage2_in_r_real_24 <= stage1_out_real_24;
stage2_in_r_imag_24  <= stage1_out_imag_24;
stage2_in_r_real_25 <= stage1_out_real_25;
stage2_in_r_imag_25  <= stage1_out_imag_25;
stage2_in_r_real_26 <= stage1_out_real_26;
stage2_in_r_imag_26  <= stage1_out_imag_26;
stage2_in_r_real_27 <= stage1_out_real_27;
stage2_in_r_imag_27  <= stage1_out_imag_27;
stage2_in_r_real_28 <= stage1_out_real_28;
stage2_in_r_imag_28  <= stage1_out_imag_28;
stage2_in_r_real_29 <= stage1_out_real_29;
stage2_in_r_imag_29  <= stage1_out_imag_29;
stage2_in_r_real_30 <= stage1_out_real_30;
stage2_in_r_imag_30  <= stage1_out_imag_30;
stage2_in_r_real_31 <= stage1_out_real_31;
stage2_in_r_imag_31  <= stage1_out_imag_31;
stage3_in_r_real_0 <= stage2_out_real_0;
stage3_in_r_imag_0  <= stage2_out_imag_0;
stage3_in_r_real_1 <= stage2_out_real_1;
stage3_in_r_imag_1  <= stage2_out_imag_1;
stage3_in_r_real_2 <= stage2_out_real_2;
stage3_in_r_imag_2  <= stage2_out_imag_2;
stage3_in_r_real_3 <= stage2_out_real_3;
stage3_in_r_imag_3  <= stage2_out_imag_3;
stage3_in_r_real_4 <= stage2_out_real_4;
stage3_in_r_imag_4  <= stage2_out_imag_4;
stage3_in_r_real_5 <= stage2_out_real_5;
stage3_in_r_imag_5  <= stage2_out_imag_5;
stage3_in_r_real_6 <= stage2_out_real_6;
stage3_in_r_imag_6  <= stage2_out_imag_6;
stage3_in_r_real_7 <= stage2_out_real_7;
stage3_in_r_imag_7  <= stage2_out_imag_7;
stage3_in_r_real_8 <= stage2_out_real_8;
stage3_in_r_imag_8  <= stage2_out_imag_8;
stage3_in_r_real_9 <= stage2_out_real_9;
stage3_in_r_imag_9  <= stage2_out_imag_9;
stage3_in_r_real_10 <= stage2_out_real_10;
stage3_in_r_imag_10  <= stage2_out_imag_10;
stage3_in_r_real_11 <= stage2_out_real_11;
stage3_in_r_imag_11  <= stage2_out_imag_11;
stage3_in_r_real_12 <= stage2_out_real_12;
stage3_in_r_imag_12  <= stage2_out_imag_12;
stage3_in_r_real_13 <= stage2_out_real_13;
stage3_in_r_imag_13  <= stage2_out_imag_13;
stage3_in_r_real_14 <= stage2_out_real_14;
stage3_in_r_imag_14  <= stage2_out_imag_14;
stage3_in_r_real_15 <= stage2_out_real_15;
stage3_in_r_imag_15  <= stage2_out_imag_15;
stage3_in_r_real_16 <= stage2_out_real_16;
stage3_in_r_imag_16  <= stage2_out_imag_16;
stage3_in_r_real_17 <= stage2_out_real_17;
stage3_in_r_imag_17  <= stage2_out_imag_17;
stage3_in_r_real_18 <= stage2_out_real_18;
stage3_in_r_imag_18  <= stage2_out_imag_18;
stage3_in_r_real_19 <= stage2_out_real_19;
stage3_in_r_imag_19  <= stage2_out_imag_19;
stage3_in_r_real_20 <= stage2_out_real_20;
stage3_in_r_imag_20  <= stage2_out_imag_20;
stage3_in_r_real_21 <= stage2_out_real_21;
stage3_in_r_imag_21  <= stage2_out_imag_21;
stage3_in_r_real_22 <= stage2_out_real_22;
stage3_in_r_imag_22  <= stage2_out_imag_22;
stage3_in_r_real_23 <= stage2_out_real_23;
stage3_in_r_imag_23  <= stage2_out_imag_23;
stage3_in_r_real_24 <= stage2_out_real_24;
stage3_in_r_imag_24  <= stage2_out_imag_24;
stage3_in_r_real_25 <= stage2_out_real_25;
stage3_in_r_imag_25  <= stage2_out_imag_25;
stage3_in_r_real_26 <= stage2_out_real_26;
stage3_in_r_imag_26  <= stage2_out_imag_26;
stage3_in_r_real_27 <= stage2_out_real_27;
stage3_in_r_imag_27  <= stage2_out_imag_27;
stage3_in_r_real_28 <= stage2_out_real_28;
stage3_in_r_imag_28  <= stage2_out_imag_28;
stage3_in_r_real_29 <= stage2_out_real_29;
stage3_in_r_imag_29  <= stage2_out_imag_29;
stage3_in_r_real_30 <= stage2_out_real_30;
stage3_in_r_imag_30  <= stage2_out_imag_30;
stage3_in_r_real_31 <= stage2_out_real_31;
stage3_in_r_imag_31  <= stage2_out_imag_31;
stage4_in_r_real_0 <= stage3_out_real_0;
stage4_in_r_imag_0  <= stage3_out_imag_0;
stage4_in_r_real_1 <= stage3_out_real_1;
stage4_in_r_imag_1  <= stage3_out_imag_1;
stage4_in_r_real_2 <= stage3_out_real_2;
stage4_in_r_imag_2  <= stage3_out_imag_2;
stage4_in_r_real_3 <= stage3_out_real_3;
stage4_in_r_imag_3  <= stage3_out_imag_3;
stage4_in_r_real_4 <= stage3_out_real_4;
stage4_in_r_imag_4  <= stage3_out_imag_4;
stage4_in_r_real_5 <= stage3_out_real_5;
stage4_in_r_imag_5  <= stage3_out_imag_5;
stage4_in_r_real_6 <= stage3_out_real_6;
stage4_in_r_imag_6  <= stage3_out_imag_6;
stage4_in_r_real_7 <= stage3_out_real_7;
stage4_in_r_imag_7  <= stage3_out_imag_7;
stage4_in_r_real_8 <= stage3_out_real_8;
stage4_in_r_imag_8  <= stage3_out_imag_8;
stage4_in_r_real_9 <= stage3_out_real_9;
stage4_in_r_imag_9  <= stage3_out_imag_9;
stage4_in_r_real_10 <= stage3_out_real_10;
stage4_in_r_imag_10  <= stage3_out_imag_10;
stage4_in_r_real_11 <= stage3_out_real_11;
stage4_in_r_imag_11  <= stage3_out_imag_11;
stage4_in_r_real_12 <= stage3_out_real_12;
stage4_in_r_imag_12  <= stage3_out_imag_12;
stage4_in_r_real_13 <= stage3_out_real_13;
stage4_in_r_imag_13  <= stage3_out_imag_13;
stage4_in_r_real_14 <= stage3_out_real_14;
stage4_in_r_imag_14  <= stage3_out_imag_14;
stage4_in_r_real_15 <= stage3_out_real_15;
stage4_in_r_imag_15  <= stage3_out_imag_15;
stage4_in_r_real_16 <= stage3_out_real_16;
stage4_in_r_imag_16  <= stage3_out_imag_16;
stage4_in_r_real_17 <= stage3_out_real_17;
stage4_in_r_imag_17  <= stage3_out_imag_17;
stage4_in_r_real_18 <= stage3_out_real_18;
stage4_in_r_imag_18  <= stage3_out_imag_18;
stage4_in_r_real_19 <= stage3_out_real_19;
stage4_in_r_imag_19  <= stage3_out_imag_19;
stage4_in_r_real_20 <= stage3_out_real_20;
stage4_in_r_imag_20  <= stage3_out_imag_20;
stage4_in_r_real_21 <= stage3_out_real_21;
stage4_in_r_imag_21  <= stage3_out_imag_21;
stage4_in_r_real_22 <= stage3_out_real_22;
stage4_in_r_imag_22  <= stage3_out_imag_22;
stage4_in_r_real_23 <= stage3_out_real_23;
stage4_in_r_imag_23  <= stage3_out_imag_23;
stage4_in_r_real_24 <= stage3_out_real_24;
stage4_in_r_imag_24  <= stage3_out_imag_24;
stage4_in_r_real_25 <= stage3_out_real_25;
stage4_in_r_imag_25  <= stage3_out_imag_25;
stage4_in_r_real_26 <= stage3_out_real_26;
stage4_in_r_imag_26  <= stage3_out_imag_26;
stage4_in_r_real_27 <= stage3_out_real_27;
stage4_in_r_imag_27  <= stage3_out_imag_27;
stage4_in_r_real_28 <= stage3_out_real_28;
stage4_in_r_imag_28  <= stage3_out_imag_28;
stage4_in_r_real_29 <= stage3_out_real_29;
stage4_in_r_imag_29  <= stage3_out_imag_29;
stage4_in_r_real_30 <= stage3_out_real_30;
stage4_in_r_imag_30  <= stage3_out_imag_30;
stage4_in_r_real_31 <= stage3_out_real_31;
stage4_in_r_imag_31  <= stage3_out_imag_31;



stage5_in_r_real_0  <= stage4_out_real_0;
stage5_in_r_imag_0 <= stage4_out_imag_0;
stage5_in_r_real_1  <= stage4_out_real_1;
stage5_in_r_imag_1 <= stage4_out_imag_1;
stage5_in_r_real_2  <= stage4_out_real_2;
stage5_in_r_imag_2 <= stage4_out_imag_2;
stage5_in_r_real_3  <= stage4_out_real_3;
stage5_in_r_imag_3 <= stage4_out_imag_3;
stage5_in_r_real_4  <= stage4_out_real_4;
stage5_in_r_imag_4 <= stage4_out_imag_4;
stage5_in_r_real_5  <= stage4_out_real_5;
stage5_in_r_imag_5 <= stage4_out_imag_5;
stage5_in_r_real_6  <= stage4_out_real_6;
stage5_in_r_imag_6 <= stage4_out_imag_6;
stage5_in_r_real_7  <= stage4_out_real_7;
stage5_in_r_imag_7 <= stage4_out_imag_7;
stage5_in_r_real_8  <= stage4_out_real_8;
stage5_in_r_imag_8 <= stage4_out_imag_8;
stage5_in_r_real_9  <= stage4_out_real_9;
stage5_in_r_imag_9 <= stage4_out_imag_9;
stage5_in_r_real_10  <= stage4_out_real_10;
stage5_in_r_imag_10 <= stage4_out_imag_10;
stage5_in_r_real_11  <= stage4_out_real_11;
stage5_in_r_imag_11 <= stage4_out_imag_11;
stage5_in_r_real_12  <= stage4_out_real_12;
stage5_in_r_imag_12 <= stage4_out_imag_12;
stage5_in_r_real_13  <= stage4_out_real_13;
stage5_in_r_imag_13 <= stage4_out_imag_13;
stage5_in_r_real_14  <= stage4_out_real_14;
stage5_in_r_imag_14 <= stage4_out_imag_14;
stage5_in_r_real_15  <= stage4_out_real_15;
stage5_in_r_imag_15 <= stage4_out_imag_15;
stage5_in_r_real_16  <= stage4_out_real_16;
stage5_in_r_imag_16 <= stage4_out_imag_16;
stage5_in_r_real_17  <= stage4_out_real_17;
stage5_in_r_imag_17 <= stage4_out_imag_17;
stage5_in_r_real_18  <= stage4_out_real_18;
stage5_in_r_imag_18 <= stage4_out_imag_18;
stage5_in_r_real_19  <= stage4_out_real_19;
stage5_in_r_imag_19 <= stage4_out_imag_19;
stage5_in_r_real_20  <= stage4_out_real_20;
stage5_in_r_imag_20 <= stage4_out_imag_20;
stage5_in_r_real_21  <= stage4_out_real_21;
stage5_in_r_imag_21 <= stage4_out_imag_21;
stage5_in_r_real_22  <= stage4_out_real_22;
stage5_in_r_imag_22 <= stage4_out_imag_22;
stage5_in_r_real_23  <= stage4_out_real_23;
stage5_in_r_imag_23 <= stage4_out_imag_23;
stage5_in_r_real_24  <= stage4_out_real_24;
stage5_in_r_imag_24 <= stage4_out_imag_24;
stage5_in_r_real_25  <= stage4_out_real_25;
stage5_in_r_imag_25 <= stage4_out_imag_25;
stage5_in_r_real_26  <= stage4_out_real_26;
stage5_in_r_imag_26 <= stage4_out_imag_26;
stage5_in_r_real_27  <= stage4_out_real_27;
stage5_in_r_imag_27 <= stage4_out_imag_27;
stage5_in_r_real_28  <= stage4_out_real_28;
stage5_in_r_imag_28 <= stage4_out_imag_28;
stage5_in_r_real_29  <= stage4_out_real_29;
stage5_in_r_imag_29 <= stage4_out_imag_29;
stage5_in_r_real_30  <= stage4_out_real_30;
stage5_in_r_imag_30 <= stage4_out_imag_30;
stage5_in_r_real_31  <= stage4_out_real_31;
stage5_in_r_imag_31 <= stage4_out_imag_31;


out_real_0 <= stage5_out_real_0;
out_imag_0 <= stage5_out_imag_0;
out_real_1 <= stage5_out_real_1;
out_imag_1 <= stage5_out_imag_1;
out_real_2 <= stage5_out_real_2;
out_imag_2 <= stage5_out_imag_2;
out_real_3 <= stage5_out_real_3;
out_imag_3 <= stage5_out_imag_3;
out_real_4 <= stage5_out_real_4;
out_imag_4 <= stage5_out_imag_4;
out_real_5 <= stage5_out_real_5;
out_imag_5 <= stage5_out_imag_5;
out_real_6 <= stage5_out_real_6;
out_imag_6 <= stage5_out_imag_6;
out_real_7 <= stage5_out_real_7;
out_imag_7 <= stage5_out_imag_7;
out_real_8 <= stage5_out_real_8;
out_imag_8 <= stage5_out_imag_8;
out_real_9 <= stage5_out_real_9;
out_imag_9 <= stage5_out_imag_9;
out_real_10 <= stage5_out_real_10;
out_imag_10 <= stage5_out_imag_10;
out_real_11 <= stage5_out_real_11;
out_imag_11 <= stage5_out_imag_11;
out_real_12 <= stage5_out_real_12;
out_imag_12 <= stage5_out_imag_12;
out_real_13 <= stage5_out_real_13;
out_imag_13 <= stage5_out_imag_13;
out_real_14 <= stage5_out_real_14;
out_imag_14 <= stage5_out_imag_14;
out_real_15 <= stage5_out_real_15;
out_imag_15 <= stage5_out_imag_15;
out_real_16 <= stage5_out_real_16;
out_imag_16 <= stage5_out_imag_16;
out_real_17 <= stage5_out_real_17;
out_imag_17 <= stage5_out_imag_17;
out_real_18 <= stage5_out_real_18;
out_imag_18 <= stage5_out_imag_18;
out_real_19 <= stage5_out_real_19;
out_imag_19 <= stage5_out_imag_19;
out_real_20 <= stage5_out_real_20;
out_imag_20 <= stage5_out_imag_20;
out_real_21 <= stage5_out_real_21;
out_imag_21 <= stage5_out_imag_21;
out_real_22 <= stage5_out_real_22;
out_imag_22 <= stage5_out_imag_22;
out_real_23 <= stage5_out_real_23;
out_imag_23 <= stage5_out_imag_23;
out_real_24 <= stage5_out_real_24;
out_imag_24 <= stage5_out_imag_24;
out_real_25 <= stage5_out_real_25;
out_imag_25 <= stage5_out_imag_25;
out_real_26 <= stage5_out_real_26;
out_imag_26 <= stage5_out_imag_26;
out_real_27 <= stage5_out_real_27;
out_imag_27 <= stage5_out_imag_27;
out_real_28 <= stage5_out_real_28;
out_imag_28 <= stage5_out_imag_28;
out_real_29 <= stage5_out_real_29;
out_imag_29 <= stage5_out_imag_29;
out_real_30 <= stage5_out_real_30;
out_imag_30 <= stage5_out_imag_30;
out_real_31 <= stage5_out_real_31;
out_imag_31 <= stage5_out_imag_31;


 end

endmodule
